`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Author: Liu Zichuan
// 
// Create Date: 09/01/2017 09:40:47 PM
// Design Name: Arthas
// Module Name: SystolicArray
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies:
// 
// Revision: 0.1
// Revision 0.01 - File Created
// Additional Comments:
//
//////////////////////////////////////////////////////////////////////////////////

module SystolicArrayWrapper(
	// inputs
	clk,
	rst,
	start,
	in_en,
	dfsm_config_en,
	dfsm_config,
	pe_config,
	pe_config_load,
	weight,
	feature,
	// outputs
	dout_en_1,
	dout_en_2,
	dout_en_3,
	dout_en_4,
	dout_en_5,
	dout_en_6,
	dout_en_7,
	dout_en_8,
	dout_en_9,
	dout_en_10,
	dout_en_11,
	dout_en_12,
	dout_en_13,
	dout_en_14,
	dout_en_15,
	dout_en_16,
	dout_en_17,
	dout_en_18,
	dout_en_19,
	dout_en_20,
	dout_en_21,
	dout_en_22,
	dout_en_23,
	dout_en_24,
	dout_en_25,
	dout_en_26,
	dout_en_27,
	dout_en_28,
	dout_en_29,
	dout_en_30,
	dout_en_31,
	dout_en_32,
	dout
);
	parameter nBanks = 11;
	parameter nCols = 32;
	parameter nRows = 3;
	parameter iWidth = 16;
	parameter oWidth = 33;
	parameter MAX_nPERIOD = 8;
	parameter MAX_nLMAC = 12288;
	parameter MAX_nSHFT = 192;

	// inputs
	input clk, rst, start, in_en, pe_config, pe_config_load, dfsm_config_en, dfsm_config;
	input [15:0] weight;
	input [15:0] feature;
	// outputs
	output dout_en_1;
	output dout_en_2;
	output dout_en_3;
	output dout_en_4;
	output dout_en_5;
	output dout_en_6;
	output dout_en_7;
	output dout_en_8;
	output dout_en_9;
	output dout_en_10;
	output dout_en_11;
	output dout_en_12;
	output dout_en_13;
	output dout_en_14;
	output dout_en_15;
	output dout_en_16;
	output dout_en_17;
	output dout_en_18;
	output dout_en_19;
	output dout_en_20;
	output dout_en_21;
	output dout_en_22;
	output dout_en_23;
	output dout_en_24;
	output dout_en_25;
	output dout_en_26;
	output dout_en_27;
	output dout_en_28;
	output dout_en_29;
	output dout_en_30;
	output dout_en_31;
	output dout_en_32;
	output [32:0] dout;

	assign dout = dout_1_1 + dout_1_2 + dout_1_3 + dout_1_4 + dout_1_5 + dout_1_6 + dout_1_7 + dout_1_8 + dout_1_9 + dout_1_10 + dout_1_11 + dout_1_12 + dout_1_13 + dout_1_14 + dout_1_15 + dout_1_16 + dout_1_17 + dout_1_18 + dout_1_19 + dout_1_20 + dout_1_21 + dout_1_22 + dout_1_23 + dout_1_24 + dout_1_25 + dout_1_26 + dout_1_27 + dout_1_28 + dout_1_29 + dout_1_30 + dout_1_31 + dout_1_32 + dout_2_1 + dout_2_2 + dout_2_3 + dout_2_4 + dout_2_5 + dout_2_6 + dout_2_7 + dout_2_8 + dout_2_9 + dout_2_10 + dout_2_11 + dout_2_12 + dout_2_13 + dout_2_14 + dout_2_15 + dout_2_16 + dout_2_17 + dout_2_18 + dout_2_19 + dout_2_20 + dout_2_21 + dout_2_22 + dout_2_23 + dout_2_24 + dout_2_25 + dout_2_26 + dout_2_27 + dout_2_28 + dout_2_29 + dout_2_30 + dout_2_31 + dout_2_32 + dout_3_1 + dout_3_2 + dout_3_3 + dout_3_4 + dout_3_5 + dout_3_6 + dout_3_7 + dout_3_8 + dout_3_9 + dout_3_10 + dout_3_11 + dout_3_12 + dout_3_13 + dout_3_14 + dout_3_15 + dout_3_16 + dout_3_17 + dout_3_18 + dout_3_19 + dout_3_20 + dout_3_21 + dout_3_22 + dout_3_23 + dout_3_24 + dout_3_25 + dout_3_26 + dout_3_27 + dout_3_28 + dout_3_29 + dout_3_30 + dout_3_31 + dout_3_32 + dout_4_1 + dout_4_2 + dout_4_3 + dout_4_4 + dout_4_5 + dout_4_6 + dout_4_7 + dout_4_8 + dout_4_9 + dout_4_10 + dout_4_11 + dout_4_12 + dout_4_13 + dout_4_14 + dout_4_15 + dout_4_16 + dout_4_17 + dout_4_18 + dout_4_19 + dout_4_20 + dout_4_21 + dout_4_22 + dout_4_23 + dout_4_24 + dout_4_25 + dout_4_26 + dout_4_27 + dout_4_28 + dout_4_29 + dout_4_30 + dout_4_31 + dout_4_32 + dout_5_1 + dout_5_2 + dout_5_3 + dout_5_4 + dout_5_5 + dout_5_6 + dout_5_7 + dout_5_8 + dout_5_9 + dout_5_10 + dout_5_11 + dout_5_12 + dout_5_13 + dout_5_14 + dout_5_15 + dout_5_16 + dout_5_17 + dout_5_18 + dout_5_19 + dout_5_20 + dout_5_21 + dout_5_22 + dout_5_23 + dout_5_24 + dout_5_25 + dout_5_26 + dout_5_27 + dout_5_28 + dout_5_29 + dout_5_30 + dout_5_31 + dout_5_32 + dout_6_1 + dout_6_2 + dout_6_3 + dout_6_4 + dout_6_5 + dout_6_6 + dout_6_7 + dout_6_8 + dout_6_9 + dout_6_10 + dout_6_11 + dout_6_12 + dout_6_13 + dout_6_14 + dout_6_15 + dout_6_16 + dout_6_17 + dout_6_18 + dout_6_19 + dout_6_20 + dout_6_21 + dout_6_22 + dout_6_23 + dout_6_24 + dout_6_25 + dout_6_26 + dout_6_27 + dout_6_28 + dout_6_29 + dout_6_30 + dout_6_31 + dout_6_32 + dout_7_1 + dout_7_2 + dout_7_3 + dout_7_4 + dout_7_5 + dout_7_6 + dout_7_7 + dout_7_8 + dout_7_9 + dout_7_10 + dout_7_11 + dout_7_12 + dout_7_13 + dout_7_14 + dout_7_15 + dout_7_16 + dout_7_17 + dout_7_18 + dout_7_19 + dout_7_20 + dout_7_21 + dout_7_22 + dout_7_23 + dout_7_24 + dout_7_25 + dout_7_26 + dout_7_27 + dout_7_28 + dout_7_29 + dout_7_30 + dout_7_31 + dout_7_32 + dout_8_1 + dout_8_2 + dout_8_3 + dout_8_4 + dout_8_5 + dout_8_6 + dout_8_7 + dout_8_8 + dout_8_9 + dout_8_10 + dout_8_11 + dout_8_12 + dout_8_13 + dout_8_14 + dout_8_15 + dout_8_16 + dout_8_17 + dout_8_18 + dout_8_19 + dout_8_20 + dout_8_21 + dout_8_22 + dout_8_23 + dout_8_24 + dout_8_25 + dout_8_26 + dout_8_27 + dout_8_28 + dout_8_29 + dout_8_30 + dout_8_31 + dout_8_32 + dout_9_1 + dout_9_2 + dout_9_3 + dout_9_4 + dout_9_5 + dout_9_6 + dout_9_7 + dout_9_8 + dout_9_9 + dout_9_10 + dout_9_11 + dout_9_12 + dout_9_13 + dout_9_14 + dout_9_15 + dout_9_16 + dout_9_17 + dout_9_18 + dout_9_19 + dout_9_20 + dout_9_21 + dout_9_22 + dout_9_23 + dout_9_24 + dout_9_25 + dout_9_26 + dout_9_27 + dout_9_28 + dout_9_29 + dout_9_30 + dout_9_31 + dout_9_32 + dout_10_1 + dout_10_2 + dout_10_3 + dout_10_4 + dout_10_5 + dout_10_6 + dout_10_7 + dout_10_8 + dout_10_9 + dout_10_10 + dout_10_11 + dout_10_12 + dout_10_13 + dout_10_14 + dout_10_15 + dout_10_16 + dout_10_17 + dout_10_18 + dout_10_19 + dout_10_20 + dout_10_21 + dout_10_22 + dout_10_23 + dout_10_24 + dout_10_25 + dout_10_26 + dout_10_27 + dout_10_28 + dout_10_29 + dout_10_30 + dout_10_31 + dout_10_32 + dout_11_1 + dout_11_2 + dout_11_3 + dout_11_4 + dout_11_5 + dout_11_6 + dout_11_7 + dout_11_8 + dout_11_9 + dout_11_10 + dout_11_11 + dout_11_12 + dout_11_13 + dout_11_14 + dout_11_15 + dout_11_16 + dout_11_17 + dout_11_18 + dout_11_19 + dout_11_20 + dout_11_21 + dout_11_22 + dout_11_23 + dout_11_24 + dout_11_25 + dout_11_26 + dout_11_27 + dout_11_28 + dout_11_29 + dout_11_30 + dout_11_31 + dout_11_32 ;

	(* KEEP = "TRUE" *) logic pe_config_1_1;
	(* KEEP = "TRUE" *) logic pe_config_1_2;
	(* KEEP = "TRUE" *) logic pe_config_1_3;
	(* KEEP = "TRUE" *) logic pe_config_2_1;
	(* KEEP = "TRUE" *) logic pe_config_2_2;
	(* KEEP = "TRUE" *) logic pe_config_2_3;
	(* KEEP = "TRUE" *) logic pe_config_3_1;
	(* KEEP = "TRUE" *) logic pe_config_3_2;
	(* KEEP = "TRUE" *) logic pe_config_3_3;
	(* KEEP = "TRUE" *) logic pe_config_4_1;
	(* KEEP = "TRUE" *) logic pe_config_4_2;
	(* KEEP = "TRUE" *) logic pe_config_4_3;
	(* KEEP = "TRUE" *) logic pe_config_5_1;
	(* KEEP = "TRUE" *) logic pe_config_5_2;
	(* KEEP = "TRUE" *) logic pe_config_5_3;
	(* KEEP = "TRUE" *) logic pe_config_6_1;
	(* KEEP = "TRUE" *) logic pe_config_6_2;
	(* KEEP = "TRUE" *) logic pe_config_6_3;
	(* KEEP = "TRUE" *) logic pe_config_7_1;
	(* KEEP = "TRUE" *) logic pe_config_7_2;
	(* KEEP = "TRUE" *) logic pe_config_7_3;
	(* KEEP = "TRUE" *) logic pe_config_8_1;
	(* KEEP = "TRUE" *) logic pe_config_8_2;
	(* KEEP = "TRUE" *) logic pe_config_8_3;
	(* KEEP = "TRUE" *) logic pe_config_9_1;
	(* KEEP = "TRUE" *) logic pe_config_9_2;
	(* KEEP = "TRUE" *) logic pe_config_9_3;
	(* KEEP = "TRUE" *) logic pe_config_10_1;
	(* KEEP = "TRUE" *) logic pe_config_10_2;
	(* KEEP = "TRUE" *) logic pe_config_10_3;
	(* KEEP = "TRUE" *) logic pe_config_11_1;
	(* KEEP = "TRUE" *) logic pe_config_11_2;
	(* KEEP = "TRUE" *) logic pe_config_11_3;
	(* KEEP = "TRUE" *) logic [15:0] weight_1_1;
	(* KEEP = "TRUE" *) logic [15:0] weight_1_2;
	(* KEEP = "TRUE" *) logic [15:0] weight_1_3;
	(* KEEP = "TRUE" *) logic [15:0] weight_2_1;
	(* KEEP = "TRUE" *) logic [15:0] weight_2_2;
	(* KEEP = "TRUE" *) logic [15:0] weight_2_3;
	(* KEEP = "TRUE" *) logic [15:0] weight_3_1;
	(* KEEP = "TRUE" *) logic [15:0] weight_3_2;
	(* KEEP = "TRUE" *) logic [15:0] weight_3_3;
	(* KEEP = "TRUE" *) logic [15:0] weight_4_1;
	(* KEEP = "TRUE" *) logic [15:0] weight_4_2;
	(* KEEP = "TRUE" *) logic [15:0] weight_4_3;
	(* KEEP = "TRUE" *) logic [15:0] weight_5_1;
	(* KEEP = "TRUE" *) logic [15:0] weight_5_2;
	(* KEEP = "TRUE" *) logic [15:0] weight_5_3;
	(* KEEP = "TRUE" *) logic [15:0] weight_6_1;
	(* KEEP = "TRUE" *) logic [15:0] weight_6_2;
	(* KEEP = "TRUE" *) logic [15:0] weight_6_3;
	(* KEEP = "TRUE" *) logic [15:0] weight_7_1;
	(* KEEP = "TRUE" *) logic [15:0] weight_7_2;
	(* KEEP = "TRUE" *) logic [15:0] weight_7_3;
	(* KEEP = "TRUE" *) logic [15:0] weight_8_1;
	(* KEEP = "TRUE" *) logic [15:0] weight_8_2;
	(* KEEP = "TRUE" *) logic [15:0] weight_8_3;
	(* KEEP = "TRUE" *) logic [15:0] weight_9_1;
	(* KEEP = "TRUE" *) logic [15:0] weight_9_2;
	(* KEEP = "TRUE" *) logic [15:0] weight_9_3;
	(* KEEP = "TRUE" *) logic [15:0] weight_10_1;
	(* KEEP = "TRUE" *) logic [15:0] weight_10_2;
	(* KEEP = "TRUE" *) logic [15:0] weight_10_3;
	(* KEEP = "TRUE" *) logic [15:0] weight_11_1;
	(* KEEP = "TRUE" *) logic [15:0] weight_11_2;
	(* KEEP = "TRUE" *) logic [15:0] weight_11_3;
	(* KEEP = "TRUE" *) logic [15:0] feature_1;
	(* KEEP = "TRUE" *) logic [15:0] feature_2;
	(* KEEP = "TRUE" *) logic [15:0] feature_3;
	(* KEEP = "TRUE" *) logic [15:0] feature_4;
	(* KEEP = "TRUE" *) logic [15:0] feature_5;
	(* KEEP = "TRUE" *) logic [15:0] feature_6;
	(* KEEP = "TRUE" *) logic [15:0] feature_7;
	(* KEEP = "TRUE" *) logic [15:0] feature_8;
	(* KEEP = "TRUE" *) logic [15:0] feature_9;
	(* KEEP = "TRUE" *) logic [15:0] feature_10;
	(* KEEP = "TRUE" *) logic [15:0] feature_11;
	(* KEEP = "TRUE" *) logic [15:0] feature_12;
	(* KEEP = "TRUE" *) logic [15:0] feature_13;
	(* KEEP = "TRUE" *) logic [15:0] feature_14;
	(* KEEP = "TRUE" *) logic [15:0] feature_15;
	(* KEEP = "TRUE" *) logic [15:0] feature_16;
	(* KEEP = "TRUE" *) logic [15:0] feature_17;
	(* KEEP = "TRUE" *) logic [15:0] feature_18;
	(* KEEP = "TRUE" *) logic [15:0] feature_19;
	(* KEEP = "TRUE" *) logic [15:0] feature_20;
	(* KEEP = "TRUE" *) logic [15:0] feature_21;
	(* KEEP = "TRUE" *) logic [15:0] feature_22;
	(* KEEP = "TRUE" *) logic [15:0] feature_23;
	(* KEEP = "TRUE" *) logic [15:0] feature_24;
	(* KEEP = "TRUE" *) logic [15:0] feature_25;
	(* KEEP = "TRUE" *) logic [15:0] feature_26;
	(* KEEP = "TRUE" *) logic [15:0] feature_27;
	(* KEEP = "TRUE" *) logic [15:0] feature_28;
	(* KEEP = "TRUE" *) logic [15:0] feature_29;
	(* KEEP = "TRUE" *) logic [15:0] feature_30;
	(* KEEP = "TRUE" *) logic [15:0] feature_31;
	(* KEEP = "TRUE" *) logic [15:0] feature_32;
	(* KEEP = "TRUE" *) logic [15:0] feature_33;
	(* KEEP = "TRUE" *) logic [15:0] feature_34;

	(* KEEP = "TRUE" *) logic [32:0] dout_1_1;
	(* KEEP = "TRUE" *) logic [32:0] dout_1_2;
	(* KEEP = "TRUE" *) logic [32:0] dout_1_3;
	(* KEEP = "TRUE" *) logic [32:0] dout_1_4;
	(* KEEP = "TRUE" *) logic [32:0] dout_1_5;
	(* KEEP = "TRUE" *) logic [32:0] dout_1_6;
	(* KEEP = "TRUE" *) logic [32:0] dout_1_7;
	(* KEEP = "TRUE" *) logic [32:0] dout_1_8;
	(* KEEP = "TRUE" *) logic [32:0] dout_1_9;
	(* KEEP = "TRUE" *) logic [32:0] dout_1_10;
	(* KEEP = "TRUE" *) logic [32:0] dout_1_11;
	(* KEEP = "TRUE" *) logic [32:0] dout_1_12;
	(* KEEP = "TRUE" *) logic [32:0] dout_1_13;
	(* KEEP = "TRUE" *) logic [32:0] dout_1_14;
	(* KEEP = "TRUE" *) logic [32:0] dout_1_15;
	(* KEEP = "TRUE" *) logic [32:0] dout_1_16;
	(* KEEP = "TRUE" *) logic [32:0] dout_1_17;
	(* KEEP = "TRUE" *) logic [32:0] dout_1_18;
	(* KEEP = "TRUE" *) logic [32:0] dout_1_19;
	(* KEEP = "TRUE" *) logic [32:0] dout_1_20;
	(* KEEP = "TRUE" *) logic [32:0] dout_1_21;
	(* KEEP = "TRUE" *) logic [32:0] dout_1_22;
	(* KEEP = "TRUE" *) logic [32:0] dout_1_23;
	(* KEEP = "TRUE" *) logic [32:0] dout_1_24;
	(* KEEP = "TRUE" *) logic [32:0] dout_1_25;
	(* KEEP = "TRUE" *) logic [32:0] dout_1_26;
	(* KEEP = "TRUE" *) logic [32:0] dout_1_27;
	(* KEEP = "TRUE" *) logic [32:0] dout_1_28;
	(* KEEP = "TRUE" *) logic [32:0] dout_1_29;
	(* KEEP = "TRUE" *) logic [32:0] dout_1_30;
	(* KEEP = "TRUE" *) logic [32:0] dout_1_31;
	(* KEEP = "TRUE" *) logic [32:0] dout_1_32;
	(* KEEP = "TRUE" *) logic [32:0] dout_2_1;
	(* KEEP = "TRUE" *) logic [32:0] dout_2_2;
	(* KEEP = "TRUE" *) logic [32:0] dout_2_3;
	(* KEEP = "TRUE" *) logic [32:0] dout_2_4;
	(* KEEP = "TRUE" *) logic [32:0] dout_2_5;
	(* KEEP = "TRUE" *) logic [32:0] dout_2_6;
	(* KEEP = "TRUE" *) logic [32:0] dout_2_7;
	(* KEEP = "TRUE" *) logic [32:0] dout_2_8;
	(* KEEP = "TRUE" *) logic [32:0] dout_2_9;
	(* KEEP = "TRUE" *) logic [32:0] dout_2_10;
	(* KEEP = "TRUE" *) logic [32:0] dout_2_11;
	(* KEEP = "TRUE" *) logic [32:0] dout_2_12;
	(* KEEP = "TRUE" *) logic [32:0] dout_2_13;
	(* KEEP = "TRUE" *) logic [32:0] dout_2_14;
	(* KEEP = "TRUE" *) logic [32:0] dout_2_15;
	(* KEEP = "TRUE" *) logic [32:0] dout_2_16;
	(* KEEP = "TRUE" *) logic [32:0] dout_2_17;
	(* KEEP = "TRUE" *) logic [32:0] dout_2_18;
	(* KEEP = "TRUE" *) logic [32:0] dout_2_19;
	(* KEEP = "TRUE" *) logic [32:0] dout_2_20;
	(* KEEP = "TRUE" *) logic [32:0] dout_2_21;
	(* KEEP = "TRUE" *) logic [32:0] dout_2_22;
	(* KEEP = "TRUE" *) logic [32:0] dout_2_23;
	(* KEEP = "TRUE" *) logic [32:0] dout_2_24;
	(* KEEP = "TRUE" *) logic [32:0] dout_2_25;
	(* KEEP = "TRUE" *) logic [32:0] dout_2_26;
	(* KEEP = "TRUE" *) logic [32:0] dout_2_27;
	(* KEEP = "TRUE" *) logic [32:0] dout_2_28;
	(* KEEP = "TRUE" *) logic [32:0] dout_2_29;
	(* KEEP = "TRUE" *) logic [32:0] dout_2_30;
	(* KEEP = "TRUE" *) logic [32:0] dout_2_31;
	(* KEEP = "TRUE" *) logic [32:0] dout_2_32;
	(* KEEP = "TRUE" *) logic [32:0] dout_3_1;
	(* KEEP = "TRUE" *) logic [32:0] dout_3_2;
	(* KEEP = "TRUE" *) logic [32:0] dout_3_3;
	(* KEEP = "TRUE" *) logic [32:0] dout_3_4;
	(* KEEP = "TRUE" *) logic [32:0] dout_3_5;
	(* KEEP = "TRUE" *) logic [32:0] dout_3_6;
	(* KEEP = "TRUE" *) logic [32:0] dout_3_7;
	(* KEEP = "TRUE" *) logic [32:0] dout_3_8;
	(* KEEP = "TRUE" *) logic [32:0] dout_3_9;
	(* KEEP = "TRUE" *) logic [32:0] dout_3_10;
	(* KEEP = "TRUE" *) logic [32:0] dout_3_11;
	(* KEEP = "TRUE" *) logic [32:0] dout_3_12;
	(* KEEP = "TRUE" *) logic [32:0] dout_3_13;
	(* KEEP = "TRUE" *) logic [32:0] dout_3_14;
	(* KEEP = "TRUE" *) logic [32:0] dout_3_15;
	(* KEEP = "TRUE" *) logic [32:0] dout_3_16;
	(* KEEP = "TRUE" *) logic [32:0] dout_3_17;
	(* KEEP = "TRUE" *) logic [32:0] dout_3_18;
	(* KEEP = "TRUE" *) logic [32:0] dout_3_19;
	(* KEEP = "TRUE" *) logic [32:0] dout_3_20;
	(* KEEP = "TRUE" *) logic [32:0] dout_3_21;
	(* KEEP = "TRUE" *) logic [32:0] dout_3_22;
	(* KEEP = "TRUE" *) logic [32:0] dout_3_23;
	(* KEEP = "TRUE" *) logic [32:0] dout_3_24;
	(* KEEP = "TRUE" *) logic [32:0] dout_3_25;
	(* KEEP = "TRUE" *) logic [32:0] dout_3_26;
	(* KEEP = "TRUE" *) logic [32:0] dout_3_27;
	(* KEEP = "TRUE" *) logic [32:0] dout_3_28;
	(* KEEP = "TRUE" *) logic [32:0] dout_3_29;
	(* KEEP = "TRUE" *) logic [32:0] dout_3_30;
	(* KEEP = "TRUE" *) logic [32:0] dout_3_31;
	(* KEEP = "TRUE" *) logic [32:0] dout_3_32;
	(* KEEP = "TRUE" *) logic [32:0] dout_4_1;
	(* KEEP = "TRUE" *) logic [32:0] dout_4_2;
	(* KEEP = "TRUE" *) logic [32:0] dout_4_3;
	(* KEEP = "TRUE" *) logic [32:0] dout_4_4;
	(* KEEP = "TRUE" *) logic [32:0] dout_4_5;
	(* KEEP = "TRUE" *) logic [32:0] dout_4_6;
	(* KEEP = "TRUE" *) logic [32:0] dout_4_7;
	(* KEEP = "TRUE" *) logic [32:0] dout_4_8;
	(* KEEP = "TRUE" *) logic [32:0] dout_4_9;
	(* KEEP = "TRUE" *) logic [32:0] dout_4_10;
	(* KEEP = "TRUE" *) logic [32:0] dout_4_11;
	(* KEEP = "TRUE" *) logic [32:0] dout_4_12;
	(* KEEP = "TRUE" *) logic [32:0] dout_4_13;
	(* KEEP = "TRUE" *) logic [32:0] dout_4_14;
	(* KEEP = "TRUE" *) logic [32:0] dout_4_15;
	(* KEEP = "TRUE" *) logic [32:0] dout_4_16;
	(* KEEP = "TRUE" *) logic [32:0] dout_4_17;
	(* KEEP = "TRUE" *) logic [32:0] dout_4_18;
	(* KEEP = "TRUE" *) logic [32:0] dout_4_19;
	(* KEEP = "TRUE" *) logic [32:0] dout_4_20;
	(* KEEP = "TRUE" *) logic [32:0] dout_4_21;
	(* KEEP = "TRUE" *) logic [32:0] dout_4_22;
	(* KEEP = "TRUE" *) logic [32:0] dout_4_23;
	(* KEEP = "TRUE" *) logic [32:0] dout_4_24;
	(* KEEP = "TRUE" *) logic [32:0] dout_4_25;
	(* KEEP = "TRUE" *) logic [32:0] dout_4_26;
	(* KEEP = "TRUE" *) logic [32:0] dout_4_27;
	(* KEEP = "TRUE" *) logic [32:0] dout_4_28;
	(* KEEP = "TRUE" *) logic [32:0] dout_4_29;
	(* KEEP = "TRUE" *) logic [32:0] dout_4_30;
	(* KEEP = "TRUE" *) logic [32:0] dout_4_31;
	(* KEEP = "TRUE" *) logic [32:0] dout_4_32;
	(* KEEP = "TRUE" *) logic [32:0] dout_5_1;
	(* KEEP = "TRUE" *) logic [32:0] dout_5_2;
	(* KEEP = "TRUE" *) logic [32:0] dout_5_3;
	(* KEEP = "TRUE" *) logic [32:0] dout_5_4;
	(* KEEP = "TRUE" *) logic [32:0] dout_5_5;
	(* KEEP = "TRUE" *) logic [32:0] dout_5_6;
	(* KEEP = "TRUE" *) logic [32:0] dout_5_7;
	(* KEEP = "TRUE" *) logic [32:0] dout_5_8;
	(* KEEP = "TRUE" *) logic [32:0] dout_5_9;
	(* KEEP = "TRUE" *) logic [32:0] dout_5_10;
	(* KEEP = "TRUE" *) logic [32:0] dout_5_11;
	(* KEEP = "TRUE" *) logic [32:0] dout_5_12;
	(* KEEP = "TRUE" *) logic [32:0] dout_5_13;
	(* KEEP = "TRUE" *) logic [32:0] dout_5_14;
	(* KEEP = "TRUE" *) logic [32:0] dout_5_15;
	(* KEEP = "TRUE" *) logic [32:0] dout_5_16;
	(* KEEP = "TRUE" *) logic [32:0] dout_5_17;
	(* KEEP = "TRUE" *) logic [32:0] dout_5_18;
	(* KEEP = "TRUE" *) logic [32:0] dout_5_19;
	(* KEEP = "TRUE" *) logic [32:0] dout_5_20;
	(* KEEP = "TRUE" *) logic [32:0] dout_5_21;
	(* KEEP = "TRUE" *) logic [32:0] dout_5_22;
	(* KEEP = "TRUE" *) logic [32:0] dout_5_23;
	(* KEEP = "TRUE" *) logic [32:0] dout_5_24;
	(* KEEP = "TRUE" *) logic [32:0] dout_5_25;
	(* KEEP = "TRUE" *) logic [32:0] dout_5_26;
	(* KEEP = "TRUE" *) logic [32:0] dout_5_27;
	(* KEEP = "TRUE" *) logic [32:0] dout_5_28;
	(* KEEP = "TRUE" *) logic [32:0] dout_5_29;
	(* KEEP = "TRUE" *) logic [32:0] dout_5_30;
	(* KEEP = "TRUE" *) logic [32:0] dout_5_31;
	(* KEEP = "TRUE" *) logic [32:0] dout_5_32;
	(* KEEP = "TRUE" *) logic [32:0] dout_6_1;
	(* KEEP = "TRUE" *) logic [32:0] dout_6_2;
	(* KEEP = "TRUE" *) logic [32:0] dout_6_3;
	(* KEEP = "TRUE" *) logic [32:0] dout_6_4;
	(* KEEP = "TRUE" *) logic [32:0] dout_6_5;
	(* KEEP = "TRUE" *) logic [32:0] dout_6_6;
	(* KEEP = "TRUE" *) logic [32:0] dout_6_7;
	(* KEEP = "TRUE" *) logic [32:0] dout_6_8;
	(* KEEP = "TRUE" *) logic [32:0] dout_6_9;
	(* KEEP = "TRUE" *) logic [32:0] dout_6_10;
	(* KEEP = "TRUE" *) logic [32:0] dout_6_11;
	(* KEEP = "TRUE" *) logic [32:0] dout_6_12;
	(* KEEP = "TRUE" *) logic [32:0] dout_6_13;
	(* KEEP = "TRUE" *) logic [32:0] dout_6_14;
	(* KEEP = "TRUE" *) logic [32:0] dout_6_15;
	(* KEEP = "TRUE" *) logic [32:0] dout_6_16;
	(* KEEP = "TRUE" *) logic [32:0] dout_6_17;
	(* KEEP = "TRUE" *) logic [32:0] dout_6_18;
	(* KEEP = "TRUE" *) logic [32:0] dout_6_19;
	(* KEEP = "TRUE" *) logic [32:0] dout_6_20;
	(* KEEP = "TRUE" *) logic [32:0] dout_6_21;
	(* KEEP = "TRUE" *) logic [32:0] dout_6_22;
	(* KEEP = "TRUE" *) logic [32:0] dout_6_23;
	(* KEEP = "TRUE" *) logic [32:0] dout_6_24;
	(* KEEP = "TRUE" *) logic [32:0] dout_6_25;
	(* KEEP = "TRUE" *) logic [32:0] dout_6_26;
	(* KEEP = "TRUE" *) logic [32:0] dout_6_27;
	(* KEEP = "TRUE" *) logic [32:0] dout_6_28;
	(* KEEP = "TRUE" *) logic [32:0] dout_6_29;
	(* KEEP = "TRUE" *) logic [32:0] dout_6_30;
	(* KEEP = "TRUE" *) logic [32:0] dout_6_31;
	(* KEEP = "TRUE" *) logic [32:0] dout_6_32;
	(* KEEP = "TRUE" *) logic [32:0] dout_7_1;
	(* KEEP = "TRUE" *) logic [32:0] dout_7_2;
	(* KEEP = "TRUE" *) logic [32:0] dout_7_3;
	(* KEEP = "TRUE" *) logic [32:0] dout_7_4;
	(* KEEP = "TRUE" *) logic [32:0] dout_7_5;
	(* KEEP = "TRUE" *) logic [32:0] dout_7_6;
	(* KEEP = "TRUE" *) logic [32:0] dout_7_7;
	(* KEEP = "TRUE" *) logic [32:0] dout_7_8;
	(* KEEP = "TRUE" *) logic [32:0] dout_7_9;
	(* KEEP = "TRUE" *) logic [32:0] dout_7_10;
	(* KEEP = "TRUE" *) logic [32:0] dout_7_11;
	(* KEEP = "TRUE" *) logic [32:0] dout_7_12;
	(* KEEP = "TRUE" *) logic [32:0] dout_7_13;
	(* KEEP = "TRUE" *) logic [32:0] dout_7_14;
	(* KEEP = "TRUE" *) logic [32:0] dout_7_15;
	(* KEEP = "TRUE" *) logic [32:0] dout_7_16;
	(* KEEP = "TRUE" *) logic [32:0] dout_7_17;
	(* KEEP = "TRUE" *) logic [32:0] dout_7_18;
	(* KEEP = "TRUE" *) logic [32:0] dout_7_19;
	(* KEEP = "TRUE" *) logic [32:0] dout_7_20;
	(* KEEP = "TRUE" *) logic [32:0] dout_7_21;
	(* KEEP = "TRUE" *) logic [32:0] dout_7_22;
	(* KEEP = "TRUE" *) logic [32:0] dout_7_23;
	(* KEEP = "TRUE" *) logic [32:0] dout_7_24;
	(* KEEP = "TRUE" *) logic [32:0] dout_7_25;
	(* KEEP = "TRUE" *) logic [32:0] dout_7_26;
	(* KEEP = "TRUE" *) logic [32:0] dout_7_27;
	(* KEEP = "TRUE" *) logic [32:0] dout_7_28;
	(* KEEP = "TRUE" *) logic [32:0] dout_7_29;
	(* KEEP = "TRUE" *) logic [32:0] dout_7_30;
	(* KEEP = "TRUE" *) logic [32:0] dout_7_31;
	(* KEEP = "TRUE" *) logic [32:0] dout_7_32;
	(* KEEP = "TRUE" *) logic [32:0] dout_8_1;
	(* KEEP = "TRUE" *) logic [32:0] dout_8_2;
	(* KEEP = "TRUE" *) logic [32:0] dout_8_3;
	(* KEEP = "TRUE" *) logic [32:0] dout_8_4;
	(* KEEP = "TRUE" *) logic [32:0] dout_8_5;
	(* KEEP = "TRUE" *) logic [32:0] dout_8_6;
	(* KEEP = "TRUE" *) logic [32:0] dout_8_7;
	(* KEEP = "TRUE" *) logic [32:0] dout_8_8;
	(* KEEP = "TRUE" *) logic [32:0] dout_8_9;
	(* KEEP = "TRUE" *) logic [32:0] dout_8_10;
	(* KEEP = "TRUE" *) logic [32:0] dout_8_11;
	(* KEEP = "TRUE" *) logic [32:0] dout_8_12;
	(* KEEP = "TRUE" *) logic [32:0] dout_8_13;
	(* KEEP = "TRUE" *) logic [32:0] dout_8_14;
	(* KEEP = "TRUE" *) logic [32:0] dout_8_15;
	(* KEEP = "TRUE" *) logic [32:0] dout_8_16;
	(* KEEP = "TRUE" *) logic [32:0] dout_8_17;
	(* KEEP = "TRUE" *) logic [32:0] dout_8_18;
	(* KEEP = "TRUE" *) logic [32:0] dout_8_19;
	(* KEEP = "TRUE" *) logic [32:0] dout_8_20;
	(* KEEP = "TRUE" *) logic [32:0] dout_8_21;
	(* KEEP = "TRUE" *) logic [32:0] dout_8_22;
	(* KEEP = "TRUE" *) logic [32:0] dout_8_23;
	(* KEEP = "TRUE" *) logic [32:0] dout_8_24;
	(* KEEP = "TRUE" *) logic [32:0] dout_8_25;
	(* KEEP = "TRUE" *) logic [32:0] dout_8_26;
	(* KEEP = "TRUE" *) logic [32:0] dout_8_27;
	(* KEEP = "TRUE" *) logic [32:0] dout_8_28;
	(* KEEP = "TRUE" *) logic [32:0] dout_8_29;
	(* KEEP = "TRUE" *) logic [32:0] dout_8_30;
	(* KEEP = "TRUE" *) logic [32:0] dout_8_31;
	(* KEEP = "TRUE" *) logic [32:0] dout_8_32;
	(* KEEP = "TRUE" *) logic [32:0] dout_9_1;
	(* KEEP = "TRUE" *) logic [32:0] dout_9_2;
	(* KEEP = "TRUE" *) logic [32:0] dout_9_3;
	(* KEEP = "TRUE" *) logic [32:0] dout_9_4;
	(* KEEP = "TRUE" *) logic [32:0] dout_9_5;
	(* KEEP = "TRUE" *) logic [32:0] dout_9_6;
	(* KEEP = "TRUE" *) logic [32:0] dout_9_7;
	(* KEEP = "TRUE" *) logic [32:0] dout_9_8;
	(* KEEP = "TRUE" *) logic [32:0] dout_9_9;
	(* KEEP = "TRUE" *) logic [32:0] dout_9_10;
	(* KEEP = "TRUE" *) logic [32:0] dout_9_11;
	(* KEEP = "TRUE" *) logic [32:0] dout_9_12;
	(* KEEP = "TRUE" *) logic [32:0] dout_9_13;
	(* KEEP = "TRUE" *) logic [32:0] dout_9_14;
	(* KEEP = "TRUE" *) logic [32:0] dout_9_15;
	(* KEEP = "TRUE" *) logic [32:0] dout_9_16;
	(* KEEP = "TRUE" *) logic [32:0] dout_9_17;
	(* KEEP = "TRUE" *) logic [32:0] dout_9_18;
	(* KEEP = "TRUE" *) logic [32:0] dout_9_19;
	(* KEEP = "TRUE" *) logic [32:0] dout_9_20;
	(* KEEP = "TRUE" *) logic [32:0] dout_9_21;
	(* KEEP = "TRUE" *) logic [32:0] dout_9_22;
	(* KEEP = "TRUE" *) logic [32:0] dout_9_23;
	(* KEEP = "TRUE" *) logic [32:0] dout_9_24;
	(* KEEP = "TRUE" *) logic [32:0] dout_9_25;
	(* KEEP = "TRUE" *) logic [32:0] dout_9_26;
	(* KEEP = "TRUE" *) logic [32:0] dout_9_27;
	(* KEEP = "TRUE" *) logic [32:0] dout_9_28;
	(* KEEP = "TRUE" *) logic [32:0] dout_9_29;
	(* KEEP = "TRUE" *) logic [32:0] dout_9_30;
	(* KEEP = "TRUE" *) logic [32:0] dout_9_31;
	(* KEEP = "TRUE" *) logic [32:0] dout_9_32;
	(* KEEP = "TRUE" *) logic [32:0] dout_10_1;
	(* KEEP = "TRUE" *) logic [32:0] dout_10_2;
	(* KEEP = "TRUE" *) logic [32:0] dout_10_3;
	(* KEEP = "TRUE" *) logic [32:0] dout_10_4;
	(* KEEP = "TRUE" *) logic [32:0] dout_10_5;
	(* KEEP = "TRUE" *) logic [32:0] dout_10_6;
	(* KEEP = "TRUE" *) logic [32:0] dout_10_7;
	(* KEEP = "TRUE" *) logic [32:0] dout_10_8;
	(* KEEP = "TRUE" *) logic [32:0] dout_10_9;
	(* KEEP = "TRUE" *) logic [32:0] dout_10_10;
	(* KEEP = "TRUE" *) logic [32:0] dout_10_11;
	(* KEEP = "TRUE" *) logic [32:0] dout_10_12;
	(* KEEP = "TRUE" *) logic [32:0] dout_10_13;
	(* KEEP = "TRUE" *) logic [32:0] dout_10_14;
	(* KEEP = "TRUE" *) logic [32:0] dout_10_15;
	(* KEEP = "TRUE" *) logic [32:0] dout_10_16;
	(* KEEP = "TRUE" *) logic [32:0] dout_10_17;
	(* KEEP = "TRUE" *) logic [32:0] dout_10_18;
	(* KEEP = "TRUE" *) logic [32:0] dout_10_19;
	(* KEEP = "TRUE" *) logic [32:0] dout_10_20;
	(* KEEP = "TRUE" *) logic [32:0] dout_10_21;
	(* KEEP = "TRUE" *) logic [32:0] dout_10_22;
	(* KEEP = "TRUE" *) logic [32:0] dout_10_23;
	(* KEEP = "TRUE" *) logic [32:0] dout_10_24;
	(* KEEP = "TRUE" *) logic [32:0] dout_10_25;
	(* KEEP = "TRUE" *) logic [32:0] dout_10_26;
	(* KEEP = "TRUE" *) logic [32:0] dout_10_27;
	(* KEEP = "TRUE" *) logic [32:0] dout_10_28;
	(* KEEP = "TRUE" *) logic [32:0] dout_10_29;
	(* KEEP = "TRUE" *) logic [32:0] dout_10_30;
	(* KEEP = "TRUE" *) logic [32:0] dout_10_31;
	(* KEEP = "TRUE" *) logic [32:0] dout_10_32;
	(* KEEP = "TRUE" *) logic [32:0] dout_11_1;
	(* KEEP = "TRUE" *) logic [32:0] dout_11_2;
	(* KEEP = "TRUE" *) logic [32:0] dout_11_3;
	(* KEEP = "TRUE" *) logic [32:0] dout_11_4;
	(* KEEP = "TRUE" *) logic [32:0] dout_11_5;
	(* KEEP = "TRUE" *) logic [32:0] dout_11_6;
	(* KEEP = "TRUE" *) logic [32:0] dout_11_7;
	(* KEEP = "TRUE" *) logic [32:0] dout_11_8;
	(* KEEP = "TRUE" *) logic [32:0] dout_11_9;
	(* KEEP = "TRUE" *) logic [32:0] dout_11_10;
	(* KEEP = "TRUE" *) logic [32:0] dout_11_11;
	(* KEEP = "TRUE" *) logic [32:0] dout_11_12;
	(* KEEP = "TRUE" *) logic [32:0] dout_11_13;
	(* KEEP = "TRUE" *) logic [32:0] dout_11_14;
	(* KEEP = "TRUE" *) logic [32:0] dout_11_15;
	(* KEEP = "TRUE" *) logic [32:0] dout_11_16;
	(* KEEP = "TRUE" *) logic [32:0] dout_11_17;
	(* KEEP = "TRUE" *) logic [32:0] dout_11_18;
	(* KEEP = "TRUE" *) logic [32:0] dout_11_19;
	(* KEEP = "TRUE" *) logic [32:0] dout_11_20;
	(* KEEP = "TRUE" *) logic [32:0] dout_11_21;
	(* KEEP = "TRUE" *) logic [32:0] dout_11_22;
	(* KEEP = "TRUE" *) logic [32:0] dout_11_23;
	(* KEEP = "TRUE" *) logic [32:0] dout_11_24;
	(* KEEP = "TRUE" *) logic [32:0] dout_11_25;
	(* KEEP = "TRUE" *) logic [32:0] dout_11_26;
	(* KEEP = "TRUE" *) logic [32:0] dout_11_27;
	(* KEEP = "TRUE" *) logic [32:0] dout_11_28;
	(* KEEP = "TRUE" *) logic [32:0] dout_11_29;
	(* KEEP = "TRUE" *) logic [32:0] dout_11_30;
	(* KEEP = "TRUE" *) logic [32:0] dout_11_31;
	(* KEEP = "TRUE" *) logic [32:0] dout_11_32;

	assign pe_config_1_1 = pe_config;
	assign pe_config_1_2 = pe_config;
	assign pe_config_1_3 = pe_config;
	assign pe_config_2_1 = pe_config;
	assign pe_config_2_2 = pe_config;
	assign pe_config_2_3 = pe_config;
	assign pe_config_3_1 = pe_config;
	assign pe_config_3_2 = pe_config;
	assign pe_config_3_3 = pe_config;
	assign pe_config_4_1 = pe_config;
	assign pe_config_4_2 = pe_config;
	assign pe_config_4_3 = pe_config;
	assign pe_config_5_1 = pe_config;
	assign pe_config_5_2 = pe_config;
	assign pe_config_5_3 = pe_config;
	assign pe_config_6_1 = pe_config;
	assign pe_config_6_2 = pe_config;
	assign pe_config_6_3 = pe_config;
	assign pe_config_7_1 = pe_config;
	assign pe_config_7_2 = pe_config;
	assign pe_config_7_3 = pe_config;
	assign pe_config_8_1 = pe_config;
	assign pe_config_8_2 = pe_config;
	assign pe_config_8_3 = pe_config;
	assign pe_config_9_1 = pe_config;
	assign pe_config_9_2 = pe_config;
	assign pe_config_9_3 = pe_config;
	assign pe_config_10_1 = pe_config;
	assign pe_config_10_2 = pe_config;
	assign pe_config_10_3 = pe_config;
	assign pe_config_11_1 = pe_config;
	assign pe_config_11_2 = pe_config;
	assign pe_config_11_3 = pe_config;

	assign weight_1_1 = weight;
	assign weight_1_2 = weight;
	assign weight_1_3 = weight;
	assign weight_2_1 = weight;
	assign weight_2_2 = weight;
	assign weight_2_3 = weight;
	assign weight_3_1 = weight;
	assign weight_3_2 = weight;
	assign weight_3_3 = weight;
	assign weight_4_1 = weight;
	assign weight_4_2 = weight;
	assign weight_4_3 = weight;
	assign weight_5_1 = weight;
	assign weight_5_2 = weight;
	assign weight_5_3 = weight;
	assign weight_6_1 = weight;
	assign weight_6_2 = weight;
	assign weight_6_3 = weight;
	assign weight_7_1 = weight;
	assign weight_7_2 = weight;
	assign weight_7_3 = weight;
	assign weight_8_1 = weight;
	assign weight_8_2 = weight;
	assign weight_8_3 = weight;
	assign weight_9_1 = weight;
	assign weight_9_2 = weight;
	assign weight_9_3 = weight;
	assign weight_10_1 = weight;
	assign weight_10_2 = weight;
	assign weight_10_3 = weight;
	assign weight_11_1 = weight;
	assign weight_11_2 = weight;
	assign weight_11_3 = weight;
	assign feature_1 = feature;
	assign feature_2 = feature;
	assign feature_3 = feature;
	assign feature_4 = feature;
	assign feature_5 = feature;
	assign feature_6 = feature;
	assign feature_7 = feature;
	assign feature_8 = feature;
	assign feature_9 = feature;
	assign feature_10 = feature;
	assign feature_11 = feature;
	assign feature_12 = feature;
	assign feature_13 = feature;
	assign feature_14 = feature;
	assign feature_15 = feature;
	assign feature_16 = feature;
	assign feature_17 = feature;
	assign feature_18 = feature;
	assign feature_19 = feature;
	assign feature_20 = feature;
	assign feature_21 = feature;
	assign feature_22 = feature;
	assign feature_23 = feature;
	assign feature_24 = feature;
	assign feature_25 = feature;
	assign feature_26 = feature;
	assign feature_27 = feature;
	assign feature_28 = feature;
	assign feature_29 = feature;
	assign feature_30 = feature;
	assign feature_31 = feature;
	assign feature_32 = feature;
	assign feature_33 = feature;
	assign feature_34 = feature;

	SystolicArray # (.iWidth(iWidth), .oWidth(oWidth), .nBanks(nBanks), .nRows(nRows), .nCols(nCols), .MAX_nPERIOD(MAX_nPERIOD), .MAX_nLMAC(MAX_nLMAC), .MAX_nSHFT(MAX_nSHFT)) U (.clk(clk), .rst(rst), .in_en(in_en), .start(start), .pe_config_1_1(pe_config_1_1), .pe_config_1_2(pe_config_1_2), .pe_config_1_3(pe_config_1_3), .pe_config_2_1(pe_config_2_1), .pe_config_2_2(pe_config_2_2), .pe_config_2_3(pe_config_2_3), .pe_config_3_1(pe_config_3_1), .pe_config_3_2(pe_config_3_2), .pe_config_3_3(pe_config_3_3), .pe_config_4_1(pe_config_4_1), .pe_config_4_2(pe_config_4_2), .pe_config_4_3(pe_config_4_3), .pe_config_5_1(pe_config_5_1), .pe_config_5_2(pe_config_5_2), .pe_config_5_3(pe_config_5_3), .pe_config_6_1(pe_config_6_1), .pe_config_6_2(pe_config_6_2), .pe_config_6_3(pe_config_6_3), .pe_config_7_1(pe_config_7_1), .pe_config_7_2(pe_config_7_2), .pe_config_7_3(pe_config_7_3), .pe_config_8_1(pe_config_8_1), .pe_config_8_2(pe_config_8_2), .pe_config_8_3(pe_config_8_3), .pe_config_9_1(pe_config_9_1), .pe_config_9_2(pe_config_9_2), .pe_config_9_3(pe_config_9_3), .pe_config_10_1(pe_config_10_1), .pe_config_10_2(pe_config_10_2), .pe_config_10_3(pe_config_10_3), .pe_config_11_1(pe_config_11_1), .pe_config_11_2(pe_config_11_2), .pe_config_11_3(pe_config_11_3), .weight_1_1(weight_1_1), .weight_1_2(weight_1_2), .weight_1_3(weight_1_3), .weight_2_1(weight_2_1), .weight_2_2(weight_2_2), .weight_2_3(weight_2_3), .weight_3_1(weight_3_1), .weight_3_2(weight_3_2), .weight_3_3(weight_3_3), .weight_4_1(weight_4_1), .weight_4_2(weight_4_2), .weight_4_3(weight_4_3), .weight_5_1(weight_5_1), .weight_5_2(weight_5_2), .weight_5_3(weight_5_3), .weight_6_1(weight_6_1), .weight_6_2(weight_6_2), .weight_6_3(weight_6_3), .weight_7_1(weight_7_1), .weight_7_2(weight_7_2), .weight_7_3(weight_7_3), .weight_8_1(weight_8_1), .weight_8_2(weight_8_2), .weight_8_3(weight_8_3), .weight_9_1(weight_9_1), .weight_9_2(weight_9_2), .weight_9_3(weight_9_3), .weight_10_1(weight_10_1), .weight_10_2(weight_10_2), .weight_10_3(weight_10_3), .weight_11_1(weight_11_1), .weight_11_2(weight_11_2), .weight_11_3(weight_11_3), .feature_1(feature_1), .feature_2(feature_2), .feature_3(feature_3), .feature_4(feature_4), .feature_5(feature_5), .feature_6(feature_6), .feature_7(feature_7), .feature_8(feature_8), .feature_9(feature_9), .feature_10(feature_10), .feature_11(feature_11), .feature_12(feature_12), .feature_13(feature_13), .feature_14(feature_14), .feature_15(feature_15), .feature_16(feature_16), .feature_17(feature_17), .feature_18(feature_18), .feature_19(feature_19), .feature_20(feature_20), .feature_21(feature_21), .feature_22(feature_22), .feature_23(feature_23), .feature_24(feature_24), .feature_25(feature_25), .feature_26(feature_26), .feature_27(feature_27), .feature_28(feature_28), .feature_29(feature_29), .feature_30(feature_30), .feature_31(feature_31), .feature_32(feature_32), .feature_33(feature_33), .feature_34(feature_34), .dout_1_1(dout_1_1), .dout_1_2(dout_1_2), .dout_1_3(dout_1_3), .dout_1_4(dout_1_4), .dout_1_5(dout_1_5), .dout_1_6(dout_1_6), .dout_1_7(dout_1_7), .dout_1_8(dout_1_8), .dout_1_9(dout_1_9), .dout_1_10(dout_1_10), .dout_1_11(dout_1_11), .dout_1_12(dout_1_12), .dout_1_13(dout_1_13), .dout_1_14(dout_1_14), .dout_1_15(dout_1_15), .dout_1_16(dout_1_16), .dout_1_17(dout_1_17), .dout_1_18(dout_1_18), .dout_1_19(dout_1_19), .dout_1_20(dout_1_20), .dout_1_21(dout_1_21), .dout_1_22(dout_1_22), .dout_1_23(dout_1_23), .dout_1_24(dout_1_24), .dout_1_25(dout_1_25), .dout_1_26(dout_1_26), .dout_1_27(dout_1_27), .dout_1_28(dout_1_28), .dout_1_29(dout_1_29), .dout_1_30(dout_1_30), .dout_1_31(dout_1_31), .dout_1_32(dout_1_32), .dout_2_1(dout_2_1), .dout_2_2(dout_2_2), .dout_2_3(dout_2_3), .dout_2_4(dout_2_4), .dout_2_5(dout_2_5), .dout_2_6(dout_2_6), .dout_2_7(dout_2_7), .dout_2_8(dout_2_8), .dout_2_9(dout_2_9), .dout_2_10(dout_2_10), .dout_2_11(dout_2_11), .dout_2_12(dout_2_12), .dout_2_13(dout_2_13), .dout_2_14(dout_2_14), .dout_2_15(dout_2_15), .dout_2_16(dout_2_16), .dout_2_17(dout_2_17), .dout_2_18(dout_2_18), .dout_2_19(dout_2_19), .dout_2_20(dout_2_20), .dout_2_21(dout_2_21), .dout_2_22(dout_2_22), .dout_2_23(dout_2_23), .dout_2_24(dout_2_24), .dout_2_25(dout_2_25), .dout_2_26(dout_2_26), .dout_2_27(dout_2_27), .dout_2_28(dout_2_28), .dout_2_29(dout_2_29), .dout_2_30(dout_2_30), .dout_2_31(dout_2_31), .dout_2_32(dout_2_32), .dout_3_1(dout_3_1), .dout_3_2(dout_3_2), .dout_3_3(dout_3_3), .dout_3_4(dout_3_4), .dout_3_5(dout_3_5), .dout_3_6(dout_3_6), .dout_3_7(dout_3_7), .dout_3_8(dout_3_8), .dout_3_9(dout_3_9), .dout_3_10(dout_3_10), .dout_3_11(dout_3_11), .dout_3_12(dout_3_12), .dout_3_13(dout_3_13), .dout_3_14(dout_3_14), .dout_3_15(dout_3_15), .dout_3_16(dout_3_16), .dout_3_17(dout_3_17), .dout_3_18(dout_3_18), .dout_3_19(dout_3_19), .dout_3_20(dout_3_20), .dout_3_21(dout_3_21), .dout_3_22(dout_3_22), .dout_3_23(dout_3_23), .dout_3_24(dout_3_24), .dout_3_25(dout_3_25), .dout_3_26(dout_3_26), .dout_3_27(dout_3_27), .dout_3_28(dout_3_28), .dout_3_29(dout_3_29), .dout_3_30(dout_3_30), .dout_3_31(dout_3_31), .dout_3_32(dout_3_32), .dout_4_1(dout_4_1), .dout_4_2(dout_4_2), .dout_4_3(dout_4_3), .dout_4_4(dout_4_4), .dout_4_5(dout_4_5), .dout_4_6(dout_4_6), .dout_4_7(dout_4_7), .dout_4_8(dout_4_8), .dout_4_9(dout_4_9), .dout_4_10(dout_4_10), .dout_4_11(dout_4_11), .dout_4_12(dout_4_12), .dout_4_13(dout_4_13), .dout_4_14(dout_4_14), .dout_4_15(dout_4_15), .dout_4_16(dout_4_16), .dout_4_17(dout_4_17), .dout_4_18(dout_4_18), .dout_4_19(dout_4_19), .dout_4_20(dout_4_20), .dout_4_21(dout_4_21), .dout_4_22(dout_4_22), .dout_4_23(dout_4_23), .dout_4_24(dout_4_24), .dout_4_25(dout_4_25), .dout_4_26(dout_4_26), .dout_4_27(dout_4_27), .dout_4_28(dout_4_28), .dout_4_29(dout_4_29), .dout_4_30(dout_4_30), .dout_4_31(dout_4_31), .dout_4_32(dout_4_32), .dout_5_1(dout_5_1), .dout_5_2(dout_5_2), .dout_5_3(dout_5_3), .dout_5_4(dout_5_4), .dout_5_5(dout_5_5), .dout_5_6(dout_5_6), .dout_5_7(dout_5_7), .dout_5_8(dout_5_8), .dout_5_9(dout_5_9), .dout_5_10(dout_5_10), .dout_5_11(dout_5_11), .dout_5_12(dout_5_12), .dout_5_13(dout_5_13), .dout_5_14(dout_5_14), .dout_5_15(dout_5_15), .dout_5_16(dout_5_16), .dout_5_17(dout_5_17), .dout_5_18(dout_5_18), .dout_5_19(dout_5_19), .dout_5_20(dout_5_20), .dout_5_21(dout_5_21), .dout_5_22(dout_5_22), .dout_5_23(dout_5_23), .dout_5_24(dout_5_24), .dout_5_25(dout_5_25), .dout_5_26(dout_5_26), .dout_5_27(dout_5_27), .dout_5_28(dout_5_28), .dout_5_29(dout_5_29), .dout_5_30(dout_5_30), .dout_5_31(dout_5_31), .dout_5_32(dout_5_32), .dout_6_1(dout_6_1), .dout_6_2(dout_6_2), .dout_6_3(dout_6_3), .dout_6_4(dout_6_4), .dout_6_5(dout_6_5), .dout_6_6(dout_6_6), .dout_6_7(dout_6_7), .dout_6_8(dout_6_8), .dout_6_9(dout_6_9), .dout_6_10(dout_6_10), .dout_6_11(dout_6_11), .dout_6_12(dout_6_12), .dout_6_13(dout_6_13), .dout_6_14(dout_6_14), .dout_6_15(dout_6_15), .dout_6_16(dout_6_16), .dout_6_17(dout_6_17), .dout_6_18(dout_6_18), .dout_6_19(dout_6_19), .dout_6_20(dout_6_20), .dout_6_21(dout_6_21), .dout_6_22(dout_6_22), .dout_6_23(dout_6_23), .dout_6_24(dout_6_24), .dout_6_25(dout_6_25), .dout_6_26(dout_6_26), .dout_6_27(dout_6_27), .dout_6_28(dout_6_28), .dout_6_29(dout_6_29), .dout_6_30(dout_6_30), .dout_6_31(dout_6_31), .dout_6_32(dout_6_32), .dout_7_1(dout_7_1), .dout_7_2(dout_7_2), .dout_7_3(dout_7_3), .dout_7_4(dout_7_4), .dout_7_5(dout_7_5), .dout_7_6(dout_7_6), .dout_7_7(dout_7_7), .dout_7_8(dout_7_8), .dout_7_9(dout_7_9), .dout_7_10(dout_7_10), .dout_7_11(dout_7_11), .dout_7_12(dout_7_12), .dout_7_13(dout_7_13), .dout_7_14(dout_7_14), .dout_7_15(dout_7_15), .dout_7_16(dout_7_16), .dout_7_17(dout_7_17), .dout_7_18(dout_7_18), .dout_7_19(dout_7_19), .dout_7_20(dout_7_20), .dout_7_21(dout_7_21), .dout_7_22(dout_7_22), .dout_7_23(dout_7_23), .dout_7_24(dout_7_24), .dout_7_25(dout_7_25), .dout_7_26(dout_7_26), .dout_7_27(dout_7_27), .dout_7_28(dout_7_28), .dout_7_29(dout_7_29), .dout_7_30(dout_7_30), .dout_7_31(dout_7_31), .dout_7_32(dout_7_32), .dout_8_1(dout_8_1), .dout_8_2(dout_8_2), .dout_8_3(dout_8_3), .dout_8_4(dout_8_4), .dout_8_5(dout_8_5), .dout_8_6(dout_8_6), .dout_8_7(dout_8_7), .dout_8_8(dout_8_8), .dout_8_9(dout_8_9), .dout_8_10(dout_8_10), .dout_8_11(dout_8_11), .dout_8_12(dout_8_12), .dout_8_13(dout_8_13), .dout_8_14(dout_8_14), .dout_8_15(dout_8_15), .dout_8_16(dout_8_16), .dout_8_17(dout_8_17), .dout_8_18(dout_8_18), .dout_8_19(dout_8_19), .dout_8_20(dout_8_20), .dout_8_21(dout_8_21), .dout_8_22(dout_8_22), .dout_8_23(dout_8_23), .dout_8_24(dout_8_24), .dout_8_25(dout_8_25), .dout_8_26(dout_8_26), .dout_8_27(dout_8_27), .dout_8_28(dout_8_28), .dout_8_29(dout_8_29), .dout_8_30(dout_8_30), .dout_8_31(dout_8_31), .dout_8_32(dout_8_32), .dout_9_1(dout_9_1), .dout_9_2(dout_9_2), .dout_9_3(dout_9_3), .dout_9_4(dout_9_4), .dout_9_5(dout_9_5), .dout_9_6(dout_9_6), .dout_9_7(dout_9_7), .dout_9_8(dout_9_8), .dout_9_9(dout_9_9), .dout_9_10(dout_9_10), .dout_9_11(dout_9_11), .dout_9_12(dout_9_12), .dout_9_13(dout_9_13), .dout_9_14(dout_9_14), .dout_9_15(dout_9_15), .dout_9_16(dout_9_16), .dout_9_17(dout_9_17), .dout_9_18(dout_9_18), .dout_9_19(dout_9_19), .dout_9_20(dout_9_20), .dout_9_21(dout_9_21), .dout_9_22(dout_9_22), .dout_9_23(dout_9_23), .dout_9_24(dout_9_24), .dout_9_25(dout_9_25), .dout_9_26(dout_9_26), .dout_9_27(dout_9_27), .dout_9_28(dout_9_28), .dout_9_29(dout_9_29), .dout_9_30(dout_9_30), .dout_9_31(dout_9_31), .dout_9_32(dout_9_32), .dout_10_1(dout_10_1), .dout_10_2(dout_10_2), .dout_10_3(dout_10_3), .dout_10_4(dout_10_4), .dout_10_5(dout_10_5), .dout_10_6(dout_10_6), .dout_10_7(dout_10_7), .dout_10_8(dout_10_8), .dout_10_9(dout_10_9), .dout_10_10(dout_10_10), .dout_10_11(dout_10_11), .dout_10_12(dout_10_12), .dout_10_13(dout_10_13), .dout_10_14(dout_10_14), .dout_10_15(dout_10_15), .dout_10_16(dout_10_16), .dout_10_17(dout_10_17), .dout_10_18(dout_10_18), .dout_10_19(dout_10_19), .dout_10_20(dout_10_20), .dout_10_21(dout_10_21), .dout_10_22(dout_10_22), .dout_10_23(dout_10_23), .dout_10_24(dout_10_24), .dout_10_25(dout_10_25), .dout_10_26(dout_10_26), .dout_10_27(dout_10_27), .dout_10_28(dout_10_28), .dout_10_29(dout_10_29), .dout_10_30(dout_10_30), .dout_10_31(dout_10_31), .dout_10_32(dout_10_32), .dout_11_1(dout_11_1), .dout_11_2(dout_11_2), .dout_11_3(dout_11_3), .dout_11_4(dout_11_4), .dout_11_5(dout_11_5), .dout_11_6(dout_11_6), .dout_11_7(dout_11_7), .dout_11_8(dout_11_8), .dout_11_9(dout_11_9), .dout_11_10(dout_11_10), .dout_11_11(dout_11_11), .dout_11_12(dout_11_12), .dout_11_13(dout_11_13), .dout_11_14(dout_11_14), .dout_11_15(dout_11_15), .dout_11_16(dout_11_16), .dout_11_17(dout_11_17), .dout_11_18(dout_11_18), .dout_11_19(dout_11_19), .dout_11_20(dout_11_20), .dout_11_21(dout_11_21), .dout_11_22(dout_11_22), .dout_11_23(dout_11_23), .dout_11_24(dout_11_24), .dout_11_25(dout_11_25), .dout_11_26(dout_11_26), .dout_11_27(dout_11_27), .dout_11_28(dout_11_28), .dout_11_29(dout_11_29), .dout_11_30(dout_11_30), .dout_11_31(dout_11_31), .dout_11_32(dout_11_32), .dout_en_1(dout_en_1), .dout_en_2(dout_en_2), .dout_en_3(dout_en_3), .dout_en_4(dout_en_4), .dout_en_5(dout_en_5), .dout_en_6(dout_en_6), .dout_en_7(dout_en_7), .dout_en_8(dout_en_8), .dout_en_9(dout_en_9), .dout_en_10(dout_en_10), .dout_en_11(dout_en_11), .dout_en_12(dout_en_12), .dout_en_13(dout_en_13), .dout_en_14(dout_en_14), .dout_en_15(dout_en_15), .dout_en_16(dout_en_16), .dout_en_17(dout_en_17), .dout_en_18(dout_en_18), .dout_en_19(dout_en_19), .dout_en_20(dout_en_20), .dout_en_21(dout_en_21), .dout_en_22(dout_en_22), .dout_en_23(dout_en_23), .dout_en_24(dout_en_24), .dout_en_25(dout_en_25), .dout_en_26(dout_en_26), .dout_en_27(dout_en_27), .dout_en_28(dout_en_28), .dout_en_29(dout_en_29), .dout_en_30(dout_en_30), .dout_en_31(dout_en_31), .dout_en_32(dout_en_32), .dfsm_config_en(dfsm_config_en), .dfsm_config(dfsm_config), .pe_config_load(pe_config_load));
endmodule
