`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: Liu Zichuan
// 
// Create Date: 09/01/2017 09:40:47 PM
// Design Name: Arthas
// Module Name: SystolicArray
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies:
// 
// Revision: 0.1
// Revision 0.01 - File Created
// Additional Comments:
//
//////////////////////////////////////////////////////////////////////////////////

module SystolicArray(
	// inputs
	clk,
	rst,
	start,
	in_en,
	dfsm_config_en,
	dfsm_config,
	pe_config_1_1,
	pe_config_1_2,
	pe_config_1_3,
	pe_config_2_1,
	pe_config_2_2,
	pe_config_2_3,
	pe_config_3_1,
	pe_config_3_2,
	pe_config_3_3,
	pe_config_4_1,
	pe_config_4_2,
	pe_config_4_3,
	pe_config_5_1,
	pe_config_5_2,
	pe_config_5_3,
	pe_config_6_1,
	pe_config_6_2,
	pe_config_6_3,
	pe_config_7_1,
	pe_config_7_2,
	pe_config_7_3,
	pe_config_8_1,
	pe_config_8_2,
	pe_config_8_3,
	pe_config_9_1,
	pe_config_9_2,
	pe_config_9_3,
	pe_config_10_1,
	pe_config_10_2,
	pe_config_10_3,
	pe_config_11_1,
	pe_config_11_2,
	pe_config_11_3,
	pe_config_load,
	weight_1_1,
	weight_1_2,
	weight_1_3,
	weight_2_1,
	weight_2_2,
	weight_2_3,
	weight_3_1,
	weight_3_2,
	weight_3_3,
	weight_4_1,
	weight_4_2,
	weight_4_3,
	weight_5_1,
	weight_5_2,
	weight_5_3,
	weight_6_1,
	weight_6_2,
	weight_6_3,
	weight_7_1,
	weight_7_2,
	weight_7_3,
	weight_8_1,
	weight_8_2,
	weight_8_3,
	weight_9_1,
	weight_9_2,
	weight_9_3,
	weight_10_1,
	weight_10_2,
	weight_10_3,
	weight_11_1,
	weight_11_2,
	weight_11_3,
	feature_1,
	feature_2,
	feature_3,
	feature_4,
	feature_5,
	feature_6,
	feature_7,
	feature_8,
	feature_9,
	feature_10,
	feature_11,
	feature_12,
	feature_13,
	feature_14,
	feature_15,
	feature_16,
	feature_17,
	feature_18,
	feature_19,
	feature_20,
	feature_21,
	feature_22,
	feature_23,
	feature_24,
	feature_25,
	feature_26,
	feature_27,
	feature_28,
	feature_29,
	feature_30,
	feature_31,
	feature_32,
	feature_33,
	feature_34,
	// outputs
	dout_1_1,
	dout_1_2,
	dout_1_3,
	dout_1_4,
	dout_1_5,
	dout_1_6,
	dout_1_7,
	dout_1_8,
	dout_1_9,
	dout_1_10,
	dout_1_11,
	dout_1_12,
	dout_1_13,
	dout_1_14,
	dout_1_15,
	dout_1_16,
	dout_1_17,
	dout_1_18,
	dout_1_19,
	dout_1_20,
	dout_1_21,
	dout_1_22,
	dout_1_23,
	dout_1_24,
	dout_1_25,
	dout_1_26,
	dout_1_27,
	dout_1_28,
	dout_1_29,
	dout_1_30,
	dout_1_31,
	dout_1_32,
	dout_2_1,
	dout_2_2,
	dout_2_3,
	dout_2_4,
	dout_2_5,
	dout_2_6,
	dout_2_7,
	dout_2_8,
	dout_2_9,
	dout_2_10,
	dout_2_11,
	dout_2_12,
	dout_2_13,
	dout_2_14,
	dout_2_15,
	dout_2_16,
	dout_2_17,
	dout_2_18,
	dout_2_19,
	dout_2_20,
	dout_2_21,
	dout_2_22,
	dout_2_23,
	dout_2_24,
	dout_2_25,
	dout_2_26,
	dout_2_27,
	dout_2_28,
	dout_2_29,
	dout_2_30,
	dout_2_31,
	dout_2_32,
	dout_3_1,
	dout_3_2,
	dout_3_3,
	dout_3_4,
	dout_3_5,
	dout_3_6,
	dout_3_7,
	dout_3_8,
	dout_3_9,
	dout_3_10,
	dout_3_11,
	dout_3_12,
	dout_3_13,
	dout_3_14,
	dout_3_15,
	dout_3_16,
	dout_3_17,
	dout_3_18,
	dout_3_19,
	dout_3_20,
	dout_3_21,
	dout_3_22,
	dout_3_23,
	dout_3_24,
	dout_3_25,
	dout_3_26,
	dout_3_27,
	dout_3_28,
	dout_3_29,
	dout_3_30,
	dout_3_31,
	dout_3_32,
	dout_4_1,
	dout_4_2,
	dout_4_3,
	dout_4_4,
	dout_4_5,
	dout_4_6,
	dout_4_7,
	dout_4_8,
	dout_4_9,
	dout_4_10,
	dout_4_11,
	dout_4_12,
	dout_4_13,
	dout_4_14,
	dout_4_15,
	dout_4_16,
	dout_4_17,
	dout_4_18,
	dout_4_19,
	dout_4_20,
	dout_4_21,
	dout_4_22,
	dout_4_23,
	dout_4_24,
	dout_4_25,
	dout_4_26,
	dout_4_27,
	dout_4_28,
	dout_4_29,
	dout_4_30,
	dout_4_31,
	dout_4_32,
	dout_5_1,
	dout_5_2,
	dout_5_3,
	dout_5_4,
	dout_5_5,
	dout_5_6,
	dout_5_7,
	dout_5_8,
	dout_5_9,
	dout_5_10,
	dout_5_11,
	dout_5_12,
	dout_5_13,
	dout_5_14,
	dout_5_15,
	dout_5_16,
	dout_5_17,
	dout_5_18,
	dout_5_19,
	dout_5_20,
	dout_5_21,
	dout_5_22,
	dout_5_23,
	dout_5_24,
	dout_5_25,
	dout_5_26,
	dout_5_27,
	dout_5_28,
	dout_5_29,
	dout_5_30,
	dout_5_31,
	dout_5_32,
	dout_6_1,
	dout_6_2,
	dout_6_3,
	dout_6_4,
	dout_6_5,
	dout_6_6,
	dout_6_7,
	dout_6_8,
	dout_6_9,
	dout_6_10,
	dout_6_11,
	dout_6_12,
	dout_6_13,
	dout_6_14,
	dout_6_15,
	dout_6_16,
	dout_6_17,
	dout_6_18,
	dout_6_19,
	dout_6_20,
	dout_6_21,
	dout_6_22,
	dout_6_23,
	dout_6_24,
	dout_6_25,
	dout_6_26,
	dout_6_27,
	dout_6_28,
	dout_6_29,
	dout_6_30,
	dout_6_31,
	dout_6_32,
	dout_7_1,
	dout_7_2,
	dout_7_3,
	dout_7_4,
	dout_7_5,
	dout_7_6,
	dout_7_7,
	dout_7_8,
	dout_7_9,
	dout_7_10,
	dout_7_11,
	dout_7_12,
	dout_7_13,
	dout_7_14,
	dout_7_15,
	dout_7_16,
	dout_7_17,
	dout_7_18,
	dout_7_19,
	dout_7_20,
	dout_7_21,
	dout_7_22,
	dout_7_23,
	dout_7_24,
	dout_7_25,
	dout_7_26,
	dout_7_27,
	dout_7_28,
	dout_7_29,
	dout_7_30,
	dout_7_31,
	dout_7_32,
	dout_8_1,
	dout_8_2,
	dout_8_3,
	dout_8_4,
	dout_8_5,
	dout_8_6,
	dout_8_7,
	dout_8_8,
	dout_8_9,
	dout_8_10,
	dout_8_11,
	dout_8_12,
	dout_8_13,
	dout_8_14,
	dout_8_15,
	dout_8_16,
	dout_8_17,
	dout_8_18,
	dout_8_19,
	dout_8_20,
	dout_8_21,
	dout_8_22,
	dout_8_23,
	dout_8_24,
	dout_8_25,
	dout_8_26,
	dout_8_27,
	dout_8_28,
	dout_8_29,
	dout_8_30,
	dout_8_31,
	dout_8_32,
	dout_9_1,
	dout_9_2,
	dout_9_3,
	dout_9_4,
	dout_9_5,
	dout_9_6,
	dout_9_7,
	dout_9_8,
	dout_9_9,
	dout_9_10,
	dout_9_11,
	dout_9_12,
	dout_9_13,
	dout_9_14,
	dout_9_15,
	dout_9_16,
	dout_9_17,
	dout_9_18,
	dout_9_19,
	dout_9_20,
	dout_9_21,
	dout_9_22,
	dout_9_23,
	dout_9_24,
	dout_9_25,
	dout_9_26,
	dout_9_27,
	dout_9_28,
	dout_9_29,
	dout_9_30,
	dout_9_31,
	dout_9_32,
	dout_10_1,
	dout_10_2,
	dout_10_3,
	dout_10_4,
	dout_10_5,
	dout_10_6,
	dout_10_7,
	dout_10_8,
	dout_10_9,
	dout_10_10,
	dout_10_11,
	dout_10_12,
	dout_10_13,
	dout_10_14,
	dout_10_15,
	dout_10_16,
	dout_10_17,
	dout_10_18,
	dout_10_19,
	dout_10_20,
	dout_10_21,
	dout_10_22,
	dout_10_23,
	dout_10_24,
	dout_10_25,
	dout_10_26,
	dout_10_27,
	dout_10_28,
	dout_10_29,
	dout_10_30,
	dout_10_31,
	dout_10_32,
	dout_11_1,
	dout_11_2,
	dout_11_3,
	dout_11_4,
	dout_11_5,
	dout_11_6,
	dout_11_7,
	dout_11_8,
	dout_11_9,
	dout_11_10,
	dout_11_11,
	dout_11_12,
	dout_11_13,
	dout_11_14,
	dout_11_15,
	dout_11_16,
	dout_11_17,
	dout_11_18,
	dout_11_19,
	dout_11_20,
	dout_11_21,
	dout_11_22,
	dout_11_23,
	dout_11_24,
	dout_11_25,
	dout_11_26,
	dout_11_27,
	dout_11_28,
	dout_11_29,
	dout_11_30,
	dout_11_31,
	dout_11_32,
	dout_en_1,
	dout_en_2,
	dout_en_3,
	dout_en_4,
	dout_en_5,
	dout_en_6,
	dout_en_7,
	dout_en_8,
	dout_en_9,
	dout_en_10,
	dout_en_11,
	dout_en_12,
	dout_en_13,
	dout_en_14,
	dout_en_15,
	dout_en_16,
	dout_en_17,
	dout_en_18,
	dout_en_19,
	dout_en_20,
	dout_en_21,
	dout_en_22,
	dout_en_23,
	dout_en_24,
	dout_en_25,
	dout_en_26,
	dout_en_27,
	dout_en_28,
	dout_en_29,
	dout_en_30,
	dout_en_31,
	dout_en_32,
);
	parameter nBanks = 11;
	parameter nCols = 32;
	parameter nRows = 3;
	parameter iWidth = 16;
	parameter oWidth = 33;
	parameter MAX_nPERIOD = 8;
	parameter MAX_nLMAC = 12288;
	parameter MAX_nSHFT = 192;

	// inputs
	input clk, rst, start, in_en, pe_config_load, dfsm_config_en, dfsm_config;
	input pe_config_1_1;
	input pe_config_1_2;
	input pe_config_1_3;
	input pe_config_2_1;
	input pe_config_2_2;
	input pe_config_2_3;
	input pe_config_3_1;
	input pe_config_3_2;
	input pe_config_3_3;
	input pe_config_4_1;
	input pe_config_4_2;
	input pe_config_4_3;
	input pe_config_5_1;
	input pe_config_5_2;
	input pe_config_5_3;
	input pe_config_6_1;
	input pe_config_6_2;
	input pe_config_6_3;
	input pe_config_7_1;
	input pe_config_7_2;
	input pe_config_7_3;
	input pe_config_8_1;
	input pe_config_8_2;
	input pe_config_8_3;
	input pe_config_9_1;
	input pe_config_9_2;
	input pe_config_9_3;
	input pe_config_10_1;
	input pe_config_10_2;
	input pe_config_10_3;
	input pe_config_11_1;
	input pe_config_11_2;
	input pe_config_11_3;
	input [15:0] weight_1_1;
	input [15:0] weight_1_2;
	input [15:0] weight_1_3;
	input [15:0] weight_2_1;
	input [15:0] weight_2_2;
	input [15:0] weight_2_3;
	input [15:0] weight_3_1;
	input [15:0] weight_3_2;
	input [15:0] weight_3_3;
	input [15:0] weight_4_1;
	input [15:0] weight_4_2;
	input [15:0] weight_4_3;
	input [15:0] weight_5_1;
	input [15:0] weight_5_2;
	input [15:0] weight_5_3;
	input [15:0] weight_6_1;
	input [15:0] weight_6_2;
	input [15:0] weight_6_3;
	input [15:0] weight_7_1;
	input [15:0] weight_7_2;
	input [15:0] weight_7_3;
	input [15:0] weight_8_1;
	input [15:0] weight_8_2;
	input [15:0] weight_8_3;
	input [15:0] weight_9_1;
	input [15:0] weight_9_2;
	input [15:0] weight_9_3;
	input [15:0] weight_10_1;
	input [15:0] weight_10_2;
	input [15:0] weight_10_3;
	input [15:0] weight_11_1;
	input [15:0] weight_11_2;
	input [15:0] weight_11_3;
	input [15:0] feature_1;
	input [15:0] feature_2;
	input [15:0] feature_3;
	input [15:0] feature_4;
	input [15:0] feature_5;
	input [15:0] feature_6;
	input [15:0] feature_7;
	input [15:0] feature_8;
	input [15:0] feature_9;
	input [15:0] feature_10;
	input [15:0] feature_11;
	input [15:0] feature_12;
	input [15:0] feature_13;
	input [15:0] feature_14;
	input [15:0] feature_15;
	input [15:0] feature_16;
	input [15:0] feature_17;
	input [15:0] feature_18;
	input [15:0] feature_19;
	input [15:0] feature_20;
	input [15:0] feature_21;
	input [15:0] feature_22;
	input [15:0] feature_23;
	input [15:0] feature_24;
	input [15:0] feature_25;
	input [15:0] feature_26;
	input [15:0] feature_27;
	input [15:0] feature_28;
	input [15:0] feature_29;
	input [15:0] feature_30;
	input [15:0] feature_31;
	input [15:0] feature_32;
	input [15:0] feature_33;
	input [15:0] feature_34;

	// outputs
	output [32:0] dout_1_1;
	output [32:0] dout_1_2;
	output [32:0] dout_1_3;
	output [32:0] dout_1_4;
	output [32:0] dout_1_5;
	output [32:0] dout_1_6;
	output [32:0] dout_1_7;
	output [32:0] dout_1_8;
	output [32:0] dout_1_9;
	output [32:0] dout_1_10;
	output [32:0] dout_1_11;
	output [32:0] dout_1_12;
	output [32:0] dout_1_13;
	output [32:0] dout_1_14;
	output [32:0] dout_1_15;
	output [32:0] dout_1_16;
	output [32:0] dout_1_17;
	output [32:0] dout_1_18;
	output [32:0] dout_1_19;
	output [32:0] dout_1_20;
	output [32:0] dout_1_21;
	output [32:0] dout_1_22;
	output [32:0] dout_1_23;
	output [32:0] dout_1_24;
	output [32:0] dout_1_25;
	output [32:0] dout_1_26;
	output [32:0] dout_1_27;
	output [32:0] dout_1_28;
	output [32:0] dout_1_29;
	output [32:0] dout_1_30;
	output [32:0] dout_1_31;
	output [32:0] dout_1_32;
	output [32:0] dout_2_1;
	output [32:0] dout_2_2;
	output [32:0] dout_2_3;
	output [32:0] dout_2_4;
	output [32:0] dout_2_5;
	output [32:0] dout_2_6;
	output [32:0] dout_2_7;
	output [32:0] dout_2_8;
	output [32:0] dout_2_9;
	output [32:0] dout_2_10;
	output [32:0] dout_2_11;
	output [32:0] dout_2_12;
	output [32:0] dout_2_13;
	output [32:0] dout_2_14;
	output [32:0] dout_2_15;
	output [32:0] dout_2_16;
	output [32:0] dout_2_17;
	output [32:0] dout_2_18;
	output [32:0] dout_2_19;
	output [32:0] dout_2_20;
	output [32:0] dout_2_21;
	output [32:0] dout_2_22;
	output [32:0] dout_2_23;
	output [32:0] dout_2_24;
	output [32:0] dout_2_25;
	output [32:0] dout_2_26;
	output [32:0] dout_2_27;
	output [32:0] dout_2_28;
	output [32:0] dout_2_29;
	output [32:0] dout_2_30;
	output [32:0] dout_2_31;
	output [32:0] dout_2_32;
	output [32:0] dout_3_1;
	output [32:0] dout_3_2;
	output [32:0] dout_3_3;
	output [32:0] dout_3_4;
	output [32:0] dout_3_5;
	output [32:0] dout_3_6;
	output [32:0] dout_3_7;
	output [32:0] dout_3_8;
	output [32:0] dout_3_9;
	output [32:0] dout_3_10;
	output [32:0] dout_3_11;
	output [32:0] dout_3_12;
	output [32:0] dout_3_13;
	output [32:0] dout_3_14;
	output [32:0] dout_3_15;
	output [32:0] dout_3_16;
	output [32:0] dout_3_17;
	output [32:0] dout_3_18;
	output [32:0] dout_3_19;
	output [32:0] dout_3_20;
	output [32:0] dout_3_21;
	output [32:0] dout_3_22;
	output [32:0] dout_3_23;
	output [32:0] dout_3_24;
	output [32:0] dout_3_25;
	output [32:0] dout_3_26;
	output [32:0] dout_3_27;
	output [32:0] dout_3_28;
	output [32:0] dout_3_29;
	output [32:0] dout_3_30;
	output [32:0] dout_3_31;
	output [32:0] dout_3_32;
	output [32:0] dout_4_1;
	output [32:0] dout_4_2;
	output [32:0] dout_4_3;
	output [32:0] dout_4_4;
	output [32:0] dout_4_5;
	output [32:0] dout_4_6;
	output [32:0] dout_4_7;
	output [32:0] dout_4_8;
	output [32:0] dout_4_9;
	output [32:0] dout_4_10;
	output [32:0] dout_4_11;
	output [32:0] dout_4_12;
	output [32:0] dout_4_13;
	output [32:0] dout_4_14;
	output [32:0] dout_4_15;
	output [32:0] dout_4_16;
	output [32:0] dout_4_17;
	output [32:0] dout_4_18;
	output [32:0] dout_4_19;
	output [32:0] dout_4_20;
	output [32:0] dout_4_21;
	output [32:0] dout_4_22;
	output [32:0] dout_4_23;
	output [32:0] dout_4_24;
	output [32:0] dout_4_25;
	output [32:0] dout_4_26;
	output [32:0] dout_4_27;
	output [32:0] dout_4_28;
	output [32:0] dout_4_29;
	output [32:0] dout_4_30;
	output [32:0] dout_4_31;
	output [32:0] dout_4_32;
	output [32:0] dout_5_1;
	output [32:0] dout_5_2;
	output [32:0] dout_5_3;
	output [32:0] dout_5_4;
	output [32:0] dout_5_5;
	output [32:0] dout_5_6;
	output [32:0] dout_5_7;
	output [32:0] dout_5_8;
	output [32:0] dout_5_9;
	output [32:0] dout_5_10;
	output [32:0] dout_5_11;
	output [32:0] dout_5_12;
	output [32:0] dout_5_13;
	output [32:0] dout_5_14;
	output [32:0] dout_5_15;
	output [32:0] dout_5_16;
	output [32:0] dout_5_17;
	output [32:0] dout_5_18;
	output [32:0] dout_5_19;
	output [32:0] dout_5_20;
	output [32:0] dout_5_21;
	output [32:0] dout_5_22;
	output [32:0] dout_5_23;
	output [32:0] dout_5_24;
	output [32:0] dout_5_25;
	output [32:0] dout_5_26;
	output [32:0] dout_5_27;
	output [32:0] dout_5_28;
	output [32:0] dout_5_29;
	output [32:0] dout_5_30;
	output [32:0] dout_5_31;
	output [32:0] dout_5_32;
	output [32:0] dout_6_1;
	output [32:0] dout_6_2;
	output [32:0] dout_6_3;
	output [32:0] dout_6_4;
	output [32:0] dout_6_5;
	output [32:0] dout_6_6;
	output [32:0] dout_6_7;
	output [32:0] dout_6_8;
	output [32:0] dout_6_9;
	output [32:0] dout_6_10;
	output [32:0] dout_6_11;
	output [32:0] dout_6_12;
	output [32:0] dout_6_13;
	output [32:0] dout_6_14;
	output [32:0] dout_6_15;
	output [32:0] dout_6_16;
	output [32:0] dout_6_17;
	output [32:0] dout_6_18;
	output [32:0] dout_6_19;
	output [32:0] dout_6_20;
	output [32:0] dout_6_21;
	output [32:0] dout_6_22;
	output [32:0] dout_6_23;
	output [32:0] dout_6_24;
	output [32:0] dout_6_25;
	output [32:0] dout_6_26;
	output [32:0] dout_6_27;
	output [32:0] dout_6_28;
	output [32:0] dout_6_29;
	output [32:0] dout_6_30;
	output [32:0] dout_6_31;
	output [32:0] dout_6_32;
	output [32:0] dout_7_1;
	output [32:0] dout_7_2;
	output [32:0] dout_7_3;
	output [32:0] dout_7_4;
	output [32:0] dout_7_5;
	output [32:0] dout_7_6;
	output [32:0] dout_7_7;
	output [32:0] dout_7_8;
	output [32:0] dout_7_9;
	output [32:0] dout_7_10;
	output [32:0] dout_7_11;
	output [32:0] dout_7_12;
	output [32:0] dout_7_13;
	output [32:0] dout_7_14;
	output [32:0] dout_7_15;
	output [32:0] dout_7_16;
	output [32:0] dout_7_17;
	output [32:0] dout_7_18;
	output [32:0] dout_7_19;
	output [32:0] dout_7_20;
	output [32:0] dout_7_21;
	output [32:0] dout_7_22;
	output [32:0] dout_7_23;
	output [32:0] dout_7_24;
	output [32:0] dout_7_25;
	output [32:0] dout_7_26;
	output [32:0] dout_7_27;
	output [32:0] dout_7_28;
	output [32:0] dout_7_29;
	output [32:0] dout_7_30;
	output [32:0] dout_7_31;
	output [32:0] dout_7_32;
	output [32:0] dout_8_1;
	output [32:0] dout_8_2;
	output [32:0] dout_8_3;
	output [32:0] dout_8_4;
	output [32:0] dout_8_5;
	output [32:0] dout_8_6;
	output [32:0] dout_8_7;
	output [32:0] dout_8_8;
	output [32:0] dout_8_9;
	output [32:0] dout_8_10;
	output [32:0] dout_8_11;
	output [32:0] dout_8_12;
	output [32:0] dout_8_13;
	output [32:0] dout_8_14;
	output [32:0] dout_8_15;
	output [32:0] dout_8_16;
	output [32:0] dout_8_17;
	output [32:0] dout_8_18;
	output [32:0] dout_8_19;
	output [32:0] dout_8_20;
	output [32:0] dout_8_21;
	output [32:0] dout_8_22;
	output [32:0] dout_8_23;
	output [32:0] dout_8_24;
	output [32:0] dout_8_25;
	output [32:0] dout_8_26;
	output [32:0] dout_8_27;
	output [32:0] dout_8_28;
	output [32:0] dout_8_29;
	output [32:0] dout_8_30;
	output [32:0] dout_8_31;
	output [32:0] dout_8_32;
	output [32:0] dout_9_1;
	output [32:0] dout_9_2;
	output [32:0] dout_9_3;
	output [32:0] dout_9_4;
	output [32:0] dout_9_5;
	output [32:0] dout_9_6;
	output [32:0] dout_9_7;
	output [32:0] dout_9_8;
	output [32:0] dout_9_9;
	output [32:0] dout_9_10;
	output [32:0] dout_9_11;
	output [32:0] dout_9_12;
	output [32:0] dout_9_13;
	output [32:0] dout_9_14;
	output [32:0] dout_9_15;
	output [32:0] dout_9_16;
	output [32:0] dout_9_17;
	output [32:0] dout_9_18;
	output [32:0] dout_9_19;
	output [32:0] dout_9_20;
	output [32:0] dout_9_21;
	output [32:0] dout_9_22;
	output [32:0] dout_9_23;
	output [32:0] dout_9_24;
	output [32:0] dout_9_25;
	output [32:0] dout_9_26;
	output [32:0] dout_9_27;
	output [32:0] dout_9_28;
	output [32:0] dout_9_29;
	output [32:0] dout_9_30;
	output [32:0] dout_9_31;
	output [32:0] dout_9_32;
	output [32:0] dout_10_1;
	output [32:0] dout_10_2;
	output [32:0] dout_10_3;
	output [32:0] dout_10_4;
	output [32:0] dout_10_5;
	output [32:0] dout_10_6;
	output [32:0] dout_10_7;
	output [32:0] dout_10_8;
	output [32:0] dout_10_9;
	output [32:0] dout_10_10;
	output [32:0] dout_10_11;
	output [32:0] dout_10_12;
	output [32:0] dout_10_13;
	output [32:0] dout_10_14;
	output [32:0] dout_10_15;
	output [32:0] dout_10_16;
	output [32:0] dout_10_17;
	output [32:0] dout_10_18;
	output [32:0] dout_10_19;
	output [32:0] dout_10_20;
	output [32:0] dout_10_21;
	output [32:0] dout_10_22;
	output [32:0] dout_10_23;
	output [32:0] dout_10_24;
	output [32:0] dout_10_25;
	output [32:0] dout_10_26;
	output [32:0] dout_10_27;
	output [32:0] dout_10_28;
	output [32:0] dout_10_29;
	output [32:0] dout_10_30;
	output [32:0] dout_10_31;
	output [32:0] dout_10_32;
	output [32:0] dout_11_1;
	output [32:0] dout_11_2;
	output [32:0] dout_11_3;
	output [32:0] dout_11_4;
	output [32:0] dout_11_5;
	output [32:0] dout_11_6;
	output [32:0] dout_11_7;
	output [32:0] dout_11_8;
	output [32:0] dout_11_9;
	output [32:0] dout_11_10;
	output [32:0] dout_11_11;
	output [32:0] dout_11_12;
	output [32:0] dout_11_13;
	output [32:0] dout_11_14;
	output [32:0] dout_11_15;
	output [32:0] dout_11_16;
	output [32:0] dout_11_17;
	output [32:0] dout_11_18;
	output [32:0] dout_11_19;
	output [32:0] dout_11_20;
	output [32:0] dout_11_21;
	output [32:0] dout_11_22;
	output [32:0] dout_11_23;
	output [32:0] dout_11_24;
	output [32:0] dout_11_25;
	output [32:0] dout_11_26;
	output [32:0] dout_11_27;
	output [32:0] dout_11_28;
	output [32:0] dout_11_29;
	output [32:0] dout_11_30;
	output [32:0] dout_11_31;
	output [32:0] dout_11_32;
	output dout_en_1;
	output dout_en_2;
	output dout_en_3;
	output dout_en_4;
	output dout_en_5;
	output dout_en_6;
	output dout_en_7;
	output dout_en_8;
	output dout_en_9;
	output dout_en_10;
	output dout_en_11;
	output dout_en_12;
	output dout_en_13;
	output dout_en_14;
	output dout_en_15;
	output dout_en_16;
	output dout_en_17;
	output dout_en_18;
	output dout_en_19;
	output dout_en_20;
	output dout_en_21;
	output dout_en_22;
	output dout_en_23;
	output dout_en_24;
	output dout_en_25;
	output dout_en_26;
	output dout_en_27;
	output dout_en_28;
	output dout_en_29;
	output dout_en_30;
	output dout_en_31;
	output dout_en_32;


	logic A_1;
	logic A_2;
	logic A_3;
	logic A_4;
	logic A_5;
	logic A_6;
	logic A_7;
	logic A_8;
	logic A_9;
	logic A_10;
	logic A_11;
	logic A_12;
	logic A_13;
	logic A_14;
	logic A_15;
	logic A_16;
	logic A_17;
	logic A_18;
	logic A_19;
	logic A_20;
	logic A_21;
	logic A_22;
	logic A_23;
	logic A_24;
	logic A_25;
	logic A_26;
	logic A_27;
	logic A_28;
	logic A_29;
	logic A_30;
	logic A_31;
	logic A_32;
	logic B_1;
	logic B_2;
	logic B_3;
	logic B_4;
	logic B_5;
	logic B_6;
	logic B_7;
	logic B_8;
	logic B_9;
	logic B_10;
	logic B_11;
	logic B_12;
	logic B_13;
	logic B_14;
	logic B_15;
	logic B_16;
	logic B_17;
	logic B_18;
	logic B_19;
	logic B_20;
	logic B_21;
	logic B_22;
	logic B_23;
	logic B_24;
	logic B_25;
	logic B_26;
	logic B_27;
	logic B_28;
	logic B_29;
	logic B_30;
	logic B_31;
	logic B_32;
	logic C_1;
	logic C_2;
	logic C_3;
	logic C_4;
	logic C_5;
	logic C_6;
	logic C_7;
	logic C_8;
	logic C_9;
	logic C_10;
	logic C_11;
	logic C_12;
	logic C_13;
	logic C_14;
	logic C_15;
	logic C_16;
	logic C_17;
	logic C_18;
	logic C_19;
	logic C_20;
	logic C_21;
	logic C_22;
	logic C_23;
	logic C_24;
	logic C_25;
	logic C_26;
	logic C_27;
	logic C_28;
	logic C_29;
	logic C_30;
	logic C_31;
	logic C_32;
	logic D_1;
	logic D_2;
	logic D_3;
	logic D_4;
	logic D_5;
	logic D_6;
	logic D_7;
	logic D_8;
	logic D_9;
	logic D_10;
	logic D_11;
	logic D_12;
	logic D_13;
	logic D_14;
	logic D_15;
	logic D_16;
	logic D_17;
	logic D_18;
	logic D_19;
	logic D_20;
	logic D_21;
	logic D_22;
	logic D_23;
	logic D_24;
	logic D_25;
	logic D_26;
	logic D_27;
	logic D_28;
	logic D_29;
	logic D_30;
	logic D_31;
	logic D_32;
	logic E_1;
	logic E_2;
	logic E_3;
	logic E_4;
	logic E_5;
	logic E_6;
	logic E_7;
	logic E_8;
	logic E_9;
	logic E_10;
	logic E_11;
	logic E_12;
	logic E_13;
	logic E_14;
	logic E_15;
	logic E_16;
	logic E_17;
	logic E_18;
	logic E_19;
	logic E_20;
	logic E_21;
	logic E_22;
	logic E_23;
	logic E_24;
	logic E_25;
	logic E_26;
	logic E_27;
	logic E_28;
	logic E_29;
	logic E_30;
	logic E_31;
	logic E_32;
	logic F_1;
	logic F_2;
	logic F_3;
	logic F_4;
	logic F_5;
	logic F_6;
	logic F_7;
	logic F_8;
	logic F_9;
	logic F_10;
	logic F_11;
	logic F_12;
	logic F_13;
	logic F_14;
	logic F_15;
	logic F_16;
	logic F_17;
	logic F_18;
	logic F_19;
	logic F_20;
	logic F_21;
	logic F_22;
	logic F_23;
	logic F_24;
	logic F_25;
	logic F_26;
	logic F_27;
	logic F_28;
	logic F_29;
	logic F_30;
	logic F_31;
	logic F_32;
	logic G_1;
	logic G_2;
	logic G_3;
	logic G_4;
	logic G_5;
	logic G_6;
	logic G_7;
	logic G_8;
	logic G_9;
	logic G_10;
	logic G_11;
	logic G_12;
	logic G_13;
	logic G_14;
	logic G_15;
	logic G_16;
	logic G_17;
	logic G_18;
	logic G_19;
	logic G_20;
	logic G_21;
	logic G_22;
	logic G_23;
	logic G_24;
	logic G_25;
	logic G_26;
	logic G_27;
	logic G_28;
	logic G_29;
	logic G_30;
	logic G_31;
	logic G_32;

	logic dfsm_data_en_1;
	logic dfsm_data_en_2;
	logic dfsm_data_en_3;
	logic dfsm_data_en_4;
	logic dfsm_data_en_5;
	logic dfsm_data_en_6;
	logic dfsm_data_en_7;
	logic dfsm_data_en_8;
	logic dfsm_data_en_9;
	logic dfsm_data_en_10;
	logic dfsm_data_en_11;
	logic dfsm_data_en_12;
	logic dfsm_data_en_13;
	logic dfsm_data_en_14;
	logic dfsm_data_en_15;
	logic dfsm_data_en_16;
	logic dfsm_data_en_17;
	logic dfsm_data_en_18;
	logic dfsm_data_en_19;
	logic dfsm_data_en_20;
	logic dfsm_data_en_21;
	logic dfsm_data_en_22;
	logic dfsm_data_en_23;
	logic dfsm_data_en_24;
	logic dfsm_data_en_25;
	logic dfsm_data_en_26;
	logic dfsm_data_en_27;
	logic dfsm_data_en_28;
	logic dfsm_data_en_29;
	logic dfsm_data_en_30;
	logic dfsm_data_en_31;
	logic dfsm_data_en_32;

	logic start_bypass_1;
	logic start_bypass_2;
	logic start_bypass_3;
	logic start_bypass_4;
	logic start_bypass_5;
	logic start_bypass_6;
	logic start_bypass_7;
	logic start_bypass_8;
	logic start_bypass_9;
	logic start_bypass_10;
	logic start_bypass_11;
	logic start_bypass_12;
	logic start_bypass_13;
	logic start_bypass_14;
	logic start_bypass_15;
	logic start_bypass_16;
	logic start_bypass_17;
	logic start_bypass_18;
	logic start_bypass_19;
	logic start_bypass_20;
	logic start_bypass_21;
	logic start_bypass_22;
	logic start_bypass_23;
	logic start_bypass_24;
	logic start_bypass_25;
	logic start_bypass_26;
	logic start_bypass_27;
	logic start_bypass_28;
	logic start_bypass_29;
	logic start_bypass_30;
	logic start_bypass_31;
	logic start_bypass_32;

	SystolicBank # (.iWidth(iWidth), .oWidth(oWidth), .nRows(nRows), .nCols(nCols)) bank_1(.clk(clk), .rst(rst), .in_en(in_en), .config_load(pe_config_load), .iconfig_1(pe_config_1_1), .iconfig_2(pe_config_1_2), .iconfig_3(pe_config_1_3), .weight_1(weight_1_1), .weight_2(weight_1_2), .weight_3(weight_1_3), .feature_1(feature_1), .feature_2(feature_2), .feature_3(feature_3), .feature_4(feature_4), .feature_5(feature_5), .feature_6(feature_6), .feature_7(feature_7), .feature_8(feature_8), .feature_9(feature_9), .feature_10(feature_10), .feature_11(feature_11), .feature_12(feature_12), .feature_13(feature_13), .feature_14(feature_14), .feature_15(feature_15), .feature_16(feature_16), .feature_17(feature_17), .feature_18(feature_18), .feature_19(feature_19), .feature_20(feature_20), .feature_21(feature_21), .feature_22(feature_22), .feature_23(feature_23), .feature_24(feature_24), .feature_25(feature_25), .feature_26(feature_26), .feature_27(feature_27), .feature_28(feature_28), .feature_29(feature_29), .feature_30(feature_30), .feature_31(feature_31), .feature_32(feature_32), .feature_33(feature_33), .feature_34(feature_34), .A_1(A_1), .A_2(A_2), .A_3(A_3), .A_4(A_4), .A_5(A_5), .A_6(A_6), .A_7(A_7), .A_8(A_8), .A_9(A_9), .A_10(A_10), .A_11(A_11), .A_12(A_12), .A_13(A_13), .A_14(A_14), .A_15(A_15), .A_16(A_16), .A_17(A_17), .A_18(A_18), .A_19(A_19), .A_20(A_20), .A_21(A_21), .A_22(A_22), .A_23(A_23), .A_24(A_24), .A_25(A_25), .A_26(A_26), .A_27(A_27), .A_28(A_28), .A_29(A_29), .A_30(A_30), .A_31(A_31), .A_32(A_32), .B_1(B_1), .B_2(B_2), .B_3(B_3), .B_4(B_4), .B_5(B_5), .B_6(B_6), .B_7(B_7), .B_8(B_8), .B_9(B_9), .B_10(B_10), .B_11(B_11), .B_12(B_12), .B_13(B_13), .B_14(B_14), .B_15(B_15), .B_16(B_16), .B_17(B_17), .B_18(B_18), .B_19(B_19), .B_20(B_20), .B_21(B_21), .B_22(B_22), .B_23(B_23), .B_24(B_24), .B_25(B_25), .B_26(B_26), .B_27(B_27), .B_28(B_28), .B_29(B_29), .B_30(B_30), .B_31(B_31), .B_32(B_32), .C_1(C_1), .C_2(C_2), .C_3(C_3), .C_4(C_4), .C_5(C_5), .C_6(C_6), .C_7(C_7), .C_8(C_8), .C_9(C_9), .C_10(C_10), .C_11(C_11), .C_12(C_12), .C_13(C_13), .C_14(C_14), .C_15(C_15), .C_16(C_16), .C_17(C_17), .C_18(C_18), .C_19(C_19), .C_20(C_20), .C_21(C_21), .C_22(C_22), .C_23(C_23), .C_24(C_24), .C_25(C_25), .C_26(C_26), .C_27(C_27), .C_28(C_28), .C_29(C_29), .C_30(C_30), .C_31(C_31), .C_32(C_32), .D_1(D_1), .D_2(D_2), .D_3(D_3), .D_4(D_4), .D_5(D_5), .D_6(D_6), .D_7(D_7), .D_8(D_8), .D_9(D_9), .D_10(D_10), .D_11(D_11), .D_12(D_12), .D_13(D_13), .D_14(D_14), .D_15(D_15), .D_16(D_16), .D_17(D_17), .D_18(D_18), .D_19(D_19), .D_20(D_20), .D_21(D_21), .D_22(D_22), .D_23(D_23), .D_24(D_24), .D_25(D_25), .D_26(D_26), .D_27(D_27), .D_28(D_28), .D_29(D_29), .D_30(D_30), .D_31(D_31), .D_32(D_32), .E_1(E_1), .E_2(E_2), .E_3(E_3), .E_4(E_4), .E_5(E_5), .E_6(E_6), .E_7(E_7), .E_8(E_8), .E_9(E_9), .E_10(E_10), .E_11(E_11), .E_12(E_12), .E_13(E_13), .E_14(E_14), .E_15(E_15), .E_16(E_16), .E_17(E_17), .E_18(E_18), .E_19(E_19), .E_20(E_20), .E_21(E_21), .E_22(E_22), .E_23(E_23), .E_24(E_24), .E_25(E_25), .E_26(E_26), .E_27(E_27), .E_28(E_28), .E_29(E_29), .E_30(E_30), .E_31(E_31), .E_32(E_32), .F_1(F_1), .F_2(F_2), .F_3(F_3), .F_4(F_4), .F_5(F_5), .F_6(F_6), .F_7(F_7), .F_8(F_8), .F_9(F_9), .F_10(F_10), .F_11(F_11), .F_12(F_12), .F_13(F_13), .F_14(F_14), .F_15(F_15), .F_16(F_16), .F_17(F_17), .F_18(F_18), .F_19(F_19), .F_20(F_20), .F_21(F_21), .F_22(F_22), .F_23(F_23), .F_24(F_24), .F_25(F_25), .F_26(F_26), .F_27(F_27), .F_28(F_28), .F_29(F_29), .F_30(F_30), .F_31(F_31), .F_32(F_32), .G_1(G_1), .G_2(G_2), .G_3(G_3), .G_4(G_4), .G_5(G_5), .G_6(G_6), .G_7(G_7), .G_8(G_8), .G_9(G_9), .G_10(G_10), .G_11(G_11), .G_12(G_12), .G_13(G_13), .G_14(G_14), .G_15(G_15), .G_16(G_16), .G_17(G_17), .G_18(G_18), .G_19(G_19), .G_20(G_20), .G_21(G_21), .G_22(G_22), .G_23(G_23), .G_24(G_24), .G_25(G_25), .G_26(G_26), .G_27(G_27), .G_28(G_28), .G_29(G_29), .G_30(G_30), .G_31(G_31), .G_32(G_32), .dout_1(dout_1_1), .dout_2(dout_1_2), .dout_3(dout_1_3), .dout_4(dout_1_4), .dout_5(dout_1_5), .dout_6(dout_1_6), .dout_7(dout_1_7), .dout_8(dout_1_8), .dout_9(dout_1_9), .dout_10(dout_1_10), .dout_11(dout_1_11), .dout_12(dout_1_12), .dout_13(dout_1_13), .dout_14(dout_1_14), .dout_15(dout_1_15), .dout_16(dout_1_16), .dout_17(dout_1_17), .dout_18(dout_1_18), .dout_19(dout_1_19), .dout_20(dout_1_20), .dout_21(dout_1_21), .dout_22(dout_1_22), .dout_23(dout_1_23), .dout_24(dout_1_24), .dout_25(dout_1_25), .dout_26(dout_1_26), .dout_27(dout_1_27), .dout_28(dout_1_28), .dout_29(dout_1_29), .dout_30(dout_1_30), .dout_31(dout_1_31), .dout_32(dout_1_32));
	SystolicBank # (.iWidth(iWidth), .oWidth(oWidth), .nRows(nRows), .nCols(nCols)) bank_2(.clk(clk), .rst(rst), .in_en(in_en), .config_load(pe_config_load), .iconfig_1(pe_config_2_1), .iconfig_2(pe_config_2_2), .iconfig_3(pe_config_2_3), .weight_1(weight_2_1), .weight_2(weight_2_2), .weight_3(weight_2_3), .feature_1(feature_1), .feature_2(feature_2), .feature_3(feature_3), .feature_4(feature_4), .feature_5(feature_5), .feature_6(feature_6), .feature_7(feature_7), .feature_8(feature_8), .feature_9(feature_9), .feature_10(feature_10), .feature_11(feature_11), .feature_12(feature_12), .feature_13(feature_13), .feature_14(feature_14), .feature_15(feature_15), .feature_16(feature_16), .feature_17(feature_17), .feature_18(feature_18), .feature_19(feature_19), .feature_20(feature_20), .feature_21(feature_21), .feature_22(feature_22), .feature_23(feature_23), .feature_24(feature_24), .feature_25(feature_25), .feature_26(feature_26), .feature_27(feature_27), .feature_28(feature_28), .feature_29(feature_29), .feature_30(feature_30), .feature_31(feature_31), .feature_32(feature_32), .feature_33(feature_33), .feature_34(feature_34), .A_1(A_1), .A_2(A_2), .A_3(A_3), .A_4(A_4), .A_5(A_5), .A_6(A_6), .A_7(A_7), .A_8(A_8), .A_9(A_9), .A_10(A_10), .A_11(A_11), .A_12(A_12), .A_13(A_13), .A_14(A_14), .A_15(A_15), .A_16(A_16), .A_17(A_17), .A_18(A_18), .A_19(A_19), .A_20(A_20), .A_21(A_21), .A_22(A_22), .A_23(A_23), .A_24(A_24), .A_25(A_25), .A_26(A_26), .A_27(A_27), .A_28(A_28), .A_29(A_29), .A_30(A_30), .A_31(A_31), .A_32(A_32), .B_1(B_1), .B_2(B_2), .B_3(B_3), .B_4(B_4), .B_5(B_5), .B_6(B_6), .B_7(B_7), .B_8(B_8), .B_9(B_9), .B_10(B_10), .B_11(B_11), .B_12(B_12), .B_13(B_13), .B_14(B_14), .B_15(B_15), .B_16(B_16), .B_17(B_17), .B_18(B_18), .B_19(B_19), .B_20(B_20), .B_21(B_21), .B_22(B_22), .B_23(B_23), .B_24(B_24), .B_25(B_25), .B_26(B_26), .B_27(B_27), .B_28(B_28), .B_29(B_29), .B_30(B_30), .B_31(B_31), .B_32(B_32), .C_1(C_1), .C_2(C_2), .C_3(C_3), .C_4(C_4), .C_5(C_5), .C_6(C_6), .C_7(C_7), .C_8(C_8), .C_9(C_9), .C_10(C_10), .C_11(C_11), .C_12(C_12), .C_13(C_13), .C_14(C_14), .C_15(C_15), .C_16(C_16), .C_17(C_17), .C_18(C_18), .C_19(C_19), .C_20(C_20), .C_21(C_21), .C_22(C_22), .C_23(C_23), .C_24(C_24), .C_25(C_25), .C_26(C_26), .C_27(C_27), .C_28(C_28), .C_29(C_29), .C_30(C_30), .C_31(C_31), .C_32(C_32), .D_1(D_1), .D_2(D_2), .D_3(D_3), .D_4(D_4), .D_5(D_5), .D_6(D_6), .D_7(D_7), .D_8(D_8), .D_9(D_9), .D_10(D_10), .D_11(D_11), .D_12(D_12), .D_13(D_13), .D_14(D_14), .D_15(D_15), .D_16(D_16), .D_17(D_17), .D_18(D_18), .D_19(D_19), .D_20(D_20), .D_21(D_21), .D_22(D_22), .D_23(D_23), .D_24(D_24), .D_25(D_25), .D_26(D_26), .D_27(D_27), .D_28(D_28), .D_29(D_29), .D_30(D_30), .D_31(D_31), .D_32(D_32), .E_1(E_1), .E_2(E_2), .E_3(E_3), .E_4(E_4), .E_5(E_5), .E_6(E_6), .E_7(E_7), .E_8(E_8), .E_9(E_9), .E_10(E_10), .E_11(E_11), .E_12(E_12), .E_13(E_13), .E_14(E_14), .E_15(E_15), .E_16(E_16), .E_17(E_17), .E_18(E_18), .E_19(E_19), .E_20(E_20), .E_21(E_21), .E_22(E_22), .E_23(E_23), .E_24(E_24), .E_25(E_25), .E_26(E_26), .E_27(E_27), .E_28(E_28), .E_29(E_29), .E_30(E_30), .E_31(E_31), .E_32(E_32), .F_1(F_1), .F_2(F_2), .F_3(F_3), .F_4(F_4), .F_5(F_5), .F_6(F_6), .F_7(F_7), .F_8(F_8), .F_9(F_9), .F_10(F_10), .F_11(F_11), .F_12(F_12), .F_13(F_13), .F_14(F_14), .F_15(F_15), .F_16(F_16), .F_17(F_17), .F_18(F_18), .F_19(F_19), .F_20(F_20), .F_21(F_21), .F_22(F_22), .F_23(F_23), .F_24(F_24), .F_25(F_25), .F_26(F_26), .F_27(F_27), .F_28(F_28), .F_29(F_29), .F_30(F_30), .F_31(F_31), .F_32(F_32), .G_1(G_1), .G_2(G_2), .G_3(G_3), .G_4(G_4), .G_5(G_5), .G_6(G_6), .G_7(G_7), .G_8(G_8), .G_9(G_9), .G_10(G_10), .G_11(G_11), .G_12(G_12), .G_13(G_13), .G_14(G_14), .G_15(G_15), .G_16(G_16), .G_17(G_17), .G_18(G_18), .G_19(G_19), .G_20(G_20), .G_21(G_21), .G_22(G_22), .G_23(G_23), .G_24(G_24), .G_25(G_25), .G_26(G_26), .G_27(G_27), .G_28(G_28), .G_29(G_29), .G_30(G_30), .G_31(G_31), .G_32(G_32), .dout_1(dout_2_1), .dout_2(dout_2_2), .dout_3(dout_2_3), .dout_4(dout_2_4), .dout_5(dout_2_5), .dout_6(dout_2_6), .dout_7(dout_2_7), .dout_8(dout_2_8), .dout_9(dout_2_9), .dout_10(dout_2_10), .dout_11(dout_2_11), .dout_12(dout_2_12), .dout_13(dout_2_13), .dout_14(dout_2_14), .dout_15(dout_2_15), .dout_16(dout_2_16), .dout_17(dout_2_17), .dout_18(dout_2_18), .dout_19(dout_2_19), .dout_20(dout_2_20), .dout_21(dout_2_21), .dout_22(dout_2_22), .dout_23(dout_2_23), .dout_24(dout_2_24), .dout_25(dout_2_25), .dout_26(dout_2_26), .dout_27(dout_2_27), .dout_28(dout_2_28), .dout_29(dout_2_29), .dout_30(dout_2_30), .dout_31(dout_2_31), .dout_32(dout_2_32));
	SystolicBank # (.iWidth(iWidth), .oWidth(oWidth), .nRows(nRows), .nCols(nCols)) bank_3(.clk(clk), .rst(rst), .in_en(in_en), .config_load(pe_config_load), .iconfig_1(pe_config_3_1), .iconfig_2(pe_config_3_2), .iconfig_3(pe_config_3_3), .weight_1(weight_3_1), .weight_2(weight_3_2), .weight_3(weight_3_3), .feature_1(feature_1), .feature_2(feature_2), .feature_3(feature_3), .feature_4(feature_4), .feature_5(feature_5), .feature_6(feature_6), .feature_7(feature_7), .feature_8(feature_8), .feature_9(feature_9), .feature_10(feature_10), .feature_11(feature_11), .feature_12(feature_12), .feature_13(feature_13), .feature_14(feature_14), .feature_15(feature_15), .feature_16(feature_16), .feature_17(feature_17), .feature_18(feature_18), .feature_19(feature_19), .feature_20(feature_20), .feature_21(feature_21), .feature_22(feature_22), .feature_23(feature_23), .feature_24(feature_24), .feature_25(feature_25), .feature_26(feature_26), .feature_27(feature_27), .feature_28(feature_28), .feature_29(feature_29), .feature_30(feature_30), .feature_31(feature_31), .feature_32(feature_32), .feature_33(feature_33), .feature_34(feature_34), .A_1(A_1), .A_2(A_2), .A_3(A_3), .A_4(A_4), .A_5(A_5), .A_6(A_6), .A_7(A_7), .A_8(A_8), .A_9(A_9), .A_10(A_10), .A_11(A_11), .A_12(A_12), .A_13(A_13), .A_14(A_14), .A_15(A_15), .A_16(A_16), .A_17(A_17), .A_18(A_18), .A_19(A_19), .A_20(A_20), .A_21(A_21), .A_22(A_22), .A_23(A_23), .A_24(A_24), .A_25(A_25), .A_26(A_26), .A_27(A_27), .A_28(A_28), .A_29(A_29), .A_30(A_30), .A_31(A_31), .A_32(A_32), .B_1(B_1), .B_2(B_2), .B_3(B_3), .B_4(B_4), .B_5(B_5), .B_6(B_6), .B_7(B_7), .B_8(B_8), .B_9(B_9), .B_10(B_10), .B_11(B_11), .B_12(B_12), .B_13(B_13), .B_14(B_14), .B_15(B_15), .B_16(B_16), .B_17(B_17), .B_18(B_18), .B_19(B_19), .B_20(B_20), .B_21(B_21), .B_22(B_22), .B_23(B_23), .B_24(B_24), .B_25(B_25), .B_26(B_26), .B_27(B_27), .B_28(B_28), .B_29(B_29), .B_30(B_30), .B_31(B_31), .B_32(B_32), .C_1(C_1), .C_2(C_2), .C_3(C_3), .C_4(C_4), .C_5(C_5), .C_6(C_6), .C_7(C_7), .C_8(C_8), .C_9(C_9), .C_10(C_10), .C_11(C_11), .C_12(C_12), .C_13(C_13), .C_14(C_14), .C_15(C_15), .C_16(C_16), .C_17(C_17), .C_18(C_18), .C_19(C_19), .C_20(C_20), .C_21(C_21), .C_22(C_22), .C_23(C_23), .C_24(C_24), .C_25(C_25), .C_26(C_26), .C_27(C_27), .C_28(C_28), .C_29(C_29), .C_30(C_30), .C_31(C_31), .C_32(C_32), .D_1(D_1), .D_2(D_2), .D_3(D_3), .D_4(D_4), .D_5(D_5), .D_6(D_6), .D_7(D_7), .D_8(D_8), .D_9(D_9), .D_10(D_10), .D_11(D_11), .D_12(D_12), .D_13(D_13), .D_14(D_14), .D_15(D_15), .D_16(D_16), .D_17(D_17), .D_18(D_18), .D_19(D_19), .D_20(D_20), .D_21(D_21), .D_22(D_22), .D_23(D_23), .D_24(D_24), .D_25(D_25), .D_26(D_26), .D_27(D_27), .D_28(D_28), .D_29(D_29), .D_30(D_30), .D_31(D_31), .D_32(D_32), .E_1(E_1), .E_2(E_2), .E_3(E_3), .E_4(E_4), .E_5(E_5), .E_6(E_6), .E_7(E_7), .E_8(E_8), .E_9(E_9), .E_10(E_10), .E_11(E_11), .E_12(E_12), .E_13(E_13), .E_14(E_14), .E_15(E_15), .E_16(E_16), .E_17(E_17), .E_18(E_18), .E_19(E_19), .E_20(E_20), .E_21(E_21), .E_22(E_22), .E_23(E_23), .E_24(E_24), .E_25(E_25), .E_26(E_26), .E_27(E_27), .E_28(E_28), .E_29(E_29), .E_30(E_30), .E_31(E_31), .E_32(E_32), .F_1(F_1), .F_2(F_2), .F_3(F_3), .F_4(F_4), .F_5(F_5), .F_6(F_6), .F_7(F_7), .F_8(F_8), .F_9(F_9), .F_10(F_10), .F_11(F_11), .F_12(F_12), .F_13(F_13), .F_14(F_14), .F_15(F_15), .F_16(F_16), .F_17(F_17), .F_18(F_18), .F_19(F_19), .F_20(F_20), .F_21(F_21), .F_22(F_22), .F_23(F_23), .F_24(F_24), .F_25(F_25), .F_26(F_26), .F_27(F_27), .F_28(F_28), .F_29(F_29), .F_30(F_30), .F_31(F_31), .F_32(F_32), .G_1(G_1), .G_2(G_2), .G_3(G_3), .G_4(G_4), .G_5(G_5), .G_6(G_6), .G_7(G_7), .G_8(G_8), .G_9(G_9), .G_10(G_10), .G_11(G_11), .G_12(G_12), .G_13(G_13), .G_14(G_14), .G_15(G_15), .G_16(G_16), .G_17(G_17), .G_18(G_18), .G_19(G_19), .G_20(G_20), .G_21(G_21), .G_22(G_22), .G_23(G_23), .G_24(G_24), .G_25(G_25), .G_26(G_26), .G_27(G_27), .G_28(G_28), .G_29(G_29), .G_30(G_30), .G_31(G_31), .G_32(G_32), .dout_1(dout_3_1), .dout_2(dout_3_2), .dout_3(dout_3_3), .dout_4(dout_3_4), .dout_5(dout_3_5), .dout_6(dout_3_6), .dout_7(dout_3_7), .dout_8(dout_3_8), .dout_9(dout_3_9), .dout_10(dout_3_10), .dout_11(dout_3_11), .dout_12(dout_3_12), .dout_13(dout_3_13), .dout_14(dout_3_14), .dout_15(dout_3_15), .dout_16(dout_3_16), .dout_17(dout_3_17), .dout_18(dout_3_18), .dout_19(dout_3_19), .dout_20(dout_3_20), .dout_21(dout_3_21), .dout_22(dout_3_22), .dout_23(dout_3_23), .dout_24(dout_3_24), .dout_25(dout_3_25), .dout_26(dout_3_26), .dout_27(dout_3_27), .dout_28(dout_3_28), .dout_29(dout_3_29), .dout_30(dout_3_30), .dout_31(dout_3_31), .dout_32(dout_3_32));
	SystolicBank # (.iWidth(iWidth), .oWidth(oWidth), .nRows(nRows), .nCols(nCols)) bank_4(.clk(clk), .rst(rst), .in_en(in_en), .config_load(pe_config_load), .iconfig_1(pe_config_4_1), .iconfig_2(pe_config_4_2), .iconfig_3(pe_config_4_3), .weight_1(weight_4_1), .weight_2(weight_4_2), .weight_3(weight_4_3), .feature_1(feature_1), .feature_2(feature_2), .feature_3(feature_3), .feature_4(feature_4), .feature_5(feature_5), .feature_6(feature_6), .feature_7(feature_7), .feature_8(feature_8), .feature_9(feature_9), .feature_10(feature_10), .feature_11(feature_11), .feature_12(feature_12), .feature_13(feature_13), .feature_14(feature_14), .feature_15(feature_15), .feature_16(feature_16), .feature_17(feature_17), .feature_18(feature_18), .feature_19(feature_19), .feature_20(feature_20), .feature_21(feature_21), .feature_22(feature_22), .feature_23(feature_23), .feature_24(feature_24), .feature_25(feature_25), .feature_26(feature_26), .feature_27(feature_27), .feature_28(feature_28), .feature_29(feature_29), .feature_30(feature_30), .feature_31(feature_31), .feature_32(feature_32), .feature_33(feature_33), .feature_34(feature_34), .A_1(A_1), .A_2(A_2), .A_3(A_3), .A_4(A_4), .A_5(A_5), .A_6(A_6), .A_7(A_7), .A_8(A_8), .A_9(A_9), .A_10(A_10), .A_11(A_11), .A_12(A_12), .A_13(A_13), .A_14(A_14), .A_15(A_15), .A_16(A_16), .A_17(A_17), .A_18(A_18), .A_19(A_19), .A_20(A_20), .A_21(A_21), .A_22(A_22), .A_23(A_23), .A_24(A_24), .A_25(A_25), .A_26(A_26), .A_27(A_27), .A_28(A_28), .A_29(A_29), .A_30(A_30), .A_31(A_31), .A_32(A_32), .B_1(B_1), .B_2(B_2), .B_3(B_3), .B_4(B_4), .B_5(B_5), .B_6(B_6), .B_7(B_7), .B_8(B_8), .B_9(B_9), .B_10(B_10), .B_11(B_11), .B_12(B_12), .B_13(B_13), .B_14(B_14), .B_15(B_15), .B_16(B_16), .B_17(B_17), .B_18(B_18), .B_19(B_19), .B_20(B_20), .B_21(B_21), .B_22(B_22), .B_23(B_23), .B_24(B_24), .B_25(B_25), .B_26(B_26), .B_27(B_27), .B_28(B_28), .B_29(B_29), .B_30(B_30), .B_31(B_31), .B_32(B_32), .C_1(C_1), .C_2(C_2), .C_3(C_3), .C_4(C_4), .C_5(C_5), .C_6(C_6), .C_7(C_7), .C_8(C_8), .C_9(C_9), .C_10(C_10), .C_11(C_11), .C_12(C_12), .C_13(C_13), .C_14(C_14), .C_15(C_15), .C_16(C_16), .C_17(C_17), .C_18(C_18), .C_19(C_19), .C_20(C_20), .C_21(C_21), .C_22(C_22), .C_23(C_23), .C_24(C_24), .C_25(C_25), .C_26(C_26), .C_27(C_27), .C_28(C_28), .C_29(C_29), .C_30(C_30), .C_31(C_31), .C_32(C_32), .D_1(D_1), .D_2(D_2), .D_3(D_3), .D_4(D_4), .D_5(D_5), .D_6(D_6), .D_7(D_7), .D_8(D_8), .D_9(D_9), .D_10(D_10), .D_11(D_11), .D_12(D_12), .D_13(D_13), .D_14(D_14), .D_15(D_15), .D_16(D_16), .D_17(D_17), .D_18(D_18), .D_19(D_19), .D_20(D_20), .D_21(D_21), .D_22(D_22), .D_23(D_23), .D_24(D_24), .D_25(D_25), .D_26(D_26), .D_27(D_27), .D_28(D_28), .D_29(D_29), .D_30(D_30), .D_31(D_31), .D_32(D_32), .E_1(E_1), .E_2(E_2), .E_3(E_3), .E_4(E_4), .E_5(E_5), .E_6(E_6), .E_7(E_7), .E_8(E_8), .E_9(E_9), .E_10(E_10), .E_11(E_11), .E_12(E_12), .E_13(E_13), .E_14(E_14), .E_15(E_15), .E_16(E_16), .E_17(E_17), .E_18(E_18), .E_19(E_19), .E_20(E_20), .E_21(E_21), .E_22(E_22), .E_23(E_23), .E_24(E_24), .E_25(E_25), .E_26(E_26), .E_27(E_27), .E_28(E_28), .E_29(E_29), .E_30(E_30), .E_31(E_31), .E_32(E_32), .F_1(F_1), .F_2(F_2), .F_3(F_3), .F_4(F_4), .F_5(F_5), .F_6(F_6), .F_7(F_7), .F_8(F_8), .F_9(F_9), .F_10(F_10), .F_11(F_11), .F_12(F_12), .F_13(F_13), .F_14(F_14), .F_15(F_15), .F_16(F_16), .F_17(F_17), .F_18(F_18), .F_19(F_19), .F_20(F_20), .F_21(F_21), .F_22(F_22), .F_23(F_23), .F_24(F_24), .F_25(F_25), .F_26(F_26), .F_27(F_27), .F_28(F_28), .F_29(F_29), .F_30(F_30), .F_31(F_31), .F_32(F_32), .G_1(G_1), .G_2(G_2), .G_3(G_3), .G_4(G_4), .G_5(G_5), .G_6(G_6), .G_7(G_7), .G_8(G_8), .G_9(G_9), .G_10(G_10), .G_11(G_11), .G_12(G_12), .G_13(G_13), .G_14(G_14), .G_15(G_15), .G_16(G_16), .G_17(G_17), .G_18(G_18), .G_19(G_19), .G_20(G_20), .G_21(G_21), .G_22(G_22), .G_23(G_23), .G_24(G_24), .G_25(G_25), .G_26(G_26), .G_27(G_27), .G_28(G_28), .G_29(G_29), .G_30(G_30), .G_31(G_31), .G_32(G_32), .dout_1(dout_4_1), .dout_2(dout_4_2), .dout_3(dout_4_3), .dout_4(dout_4_4), .dout_5(dout_4_5), .dout_6(dout_4_6), .dout_7(dout_4_7), .dout_8(dout_4_8), .dout_9(dout_4_9), .dout_10(dout_4_10), .dout_11(dout_4_11), .dout_12(dout_4_12), .dout_13(dout_4_13), .dout_14(dout_4_14), .dout_15(dout_4_15), .dout_16(dout_4_16), .dout_17(dout_4_17), .dout_18(dout_4_18), .dout_19(dout_4_19), .dout_20(dout_4_20), .dout_21(dout_4_21), .dout_22(dout_4_22), .dout_23(dout_4_23), .dout_24(dout_4_24), .dout_25(dout_4_25), .dout_26(dout_4_26), .dout_27(dout_4_27), .dout_28(dout_4_28), .dout_29(dout_4_29), .dout_30(dout_4_30), .dout_31(dout_4_31), .dout_32(dout_4_32));
	SystolicBank # (.iWidth(iWidth), .oWidth(oWidth), .nRows(nRows), .nCols(nCols)) bank_5(.clk(clk), .rst(rst), .in_en(in_en), .config_load(pe_config_load), .iconfig_1(pe_config_5_1), .iconfig_2(pe_config_5_2), .iconfig_3(pe_config_5_3), .weight_1(weight_5_1), .weight_2(weight_5_2), .weight_3(weight_5_3), .feature_1(feature_1), .feature_2(feature_2), .feature_3(feature_3), .feature_4(feature_4), .feature_5(feature_5), .feature_6(feature_6), .feature_7(feature_7), .feature_8(feature_8), .feature_9(feature_9), .feature_10(feature_10), .feature_11(feature_11), .feature_12(feature_12), .feature_13(feature_13), .feature_14(feature_14), .feature_15(feature_15), .feature_16(feature_16), .feature_17(feature_17), .feature_18(feature_18), .feature_19(feature_19), .feature_20(feature_20), .feature_21(feature_21), .feature_22(feature_22), .feature_23(feature_23), .feature_24(feature_24), .feature_25(feature_25), .feature_26(feature_26), .feature_27(feature_27), .feature_28(feature_28), .feature_29(feature_29), .feature_30(feature_30), .feature_31(feature_31), .feature_32(feature_32), .feature_33(feature_33), .feature_34(feature_34), .A_1(A_1), .A_2(A_2), .A_3(A_3), .A_4(A_4), .A_5(A_5), .A_6(A_6), .A_7(A_7), .A_8(A_8), .A_9(A_9), .A_10(A_10), .A_11(A_11), .A_12(A_12), .A_13(A_13), .A_14(A_14), .A_15(A_15), .A_16(A_16), .A_17(A_17), .A_18(A_18), .A_19(A_19), .A_20(A_20), .A_21(A_21), .A_22(A_22), .A_23(A_23), .A_24(A_24), .A_25(A_25), .A_26(A_26), .A_27(A_27), .A_28(A_28), .A_29(A_29), .A_30(A_30), .A_31(A_31), .A_32(A_32), .B_1(B_1), .B_2(B_2), .B_3(B_3), .B_4(B_4), .B_5(B_5), .B_6(B_6), .B_7(B_7), .B_8(B_8), .B_9(B_9), .B_10(B_10), .B_11(B_11), .B_12(B_12), .B_13(B_13), .B_14(B_14), .B_15(B_15), .B_16(B_16), .B_17(B_17), .B_18(B_18), .B_19(B_19), .B_20(B_20), .B_21(B_21), .B_22(B_22), .B_23(B_23), .B_24(B_24), .B_25(B_25), .B_26(B_26), .B_27(B_27), .B_28(B_28), .B_29(B_29), .B_30(B_30), .B_31(B_31), .B_32(B_32), .C_1(C_1), .C_2(C_2), .C_3(C_3), .C_4(C_4), .C_5(C_5), .C_6(C_6), .C_7(C_7), .C_8(C_8), .C_9(C_9), .C_10(C_10), .C_11(C_11), .C_12(C_12), .C_13(C_13), .C_14(C_14), .C_15(C_15), .C_16(C_16), .C_17(C_17), .C_18(C_18), .C_19(C_19), .C_20(C_20), .C_21(C_21), .C_22(C_22), .C_23(C_23), .C_24(C_24), .C_25(C_25), .C_26(C_26), .C_27(C_27), .C_28(C_28), .C_29(C_29), .C_30(C_30), .C_31(C_31), .C_32(C_32), .D_1(D_1), .D_2(D_2), .D_3(D_3), .D_4(D_4), .D_5(D_5), .D_6(D_6), .D_7(D_7), .D_8(D_8), .D_9(D_9), .D_10(D_10), .D_11(D_11), .D_12(D_12), .D_13(D_13), .D_14(D_14), .D_15(D_15), .D_16(D_16), .D_17(D_17), .D_18(D_18), .D_19(D_19), .D_20(D_20), .D_21(D_21), .D_22(D_22), .D_23(D_23), .D_24(D_24), .D_25(D_25), .D_26(D_26), .D_27(D_27), .D_28(D_28), .D_29(D_29), .D_30(D_30), .D_31(D_31), .D_32(D_32), .E_1(E_1), .E_2(E_2), .E_3(E_3), .E_4(E_4), .E_5(E_5), .E_6(E_6), .E_7(E_7), .E_8(E_8), .E_9(E_9), .E_10(E_10), .E_11(E_11), .E_12(E_12), .E_13(E_13), .E_14(E_14), .E_15(E_15), .E_16(E_16), .E_17(E_17), .E_18(E_18), .E_19(E_19), .E_20(E_20), .E_21(E_21), .E_22(E_22), .E_23(E_23), .E_24(E_24), .E_25(E_25), .E_26(E_26), .E_27(E_27), .E_28(E_28), .E_29(E_29), .E_30(E_30), .E_31(E_31), .E_32(E_32), .F_1(F_1), .F_2(F_2), .F_3(F_3), .F_4(F_4), .F_5(F_5), .F_6(F_6), .F_7(F_7), .F_8(F_8), .F_9(F_9), .F_10(F_10), .F_11(F_11), .F_12(F_12), .F_13(F_13), .F_14(F_14), .F_15(F_15), .F_16(F_16), .F_17(F_17), .F_18(F_18), .F_19(F_19), .F_20(F_20), .F_21(F_21), .F_22(F_22), .F_23(F_23), .F_24(F_24), .F_25(F_25), .F_26(F_26), .F_27(F_27), .F_28(F_28), .F_29(F_29), .F_30(F_30), .F_31(F_31), .F_32(F_32), .G_1(G_1), .G_2(G_2), .G_3(G_3), .G_4(G_4), .G_5(G_5), .G_6(G_6), .G_7(G_7), .G_8(G_8), .G_9(G_9), .G_10(G_10), .G_11(G_11), .G_12(G_12), .G_13(G_13), .G_14(G_14), .G_15(G_15), .G_16(G_16), .G_17(G_17), .G_18(G_18), .G_19(G_19), .G_20(G_20), .G_21(G_21), .G_22(G_22), .G_23(G_23), .G_24(G_24), .G_25(G_25), .G_26(G_26), .G_27(G_27), .G_28(G_28), .G_29(G_29), .G_30(G_30), .G_31(G_31), .G_32(G_32), .dout_1(dout_5_1), .dout_2(dout_5_2), .dout_3(dout_5_3), .dout_4(dout_5_4), .dout_5(dout_5_5), .dout_6(dout_5_6), .dout_7(dout_5_7), .dout_8(dout_5_8), .dout_9(dout_5_9), .dout_10(dout_5_10), .dout_11(dout_5_11), .dout_12(dout_5_12), .dout_13(dout_5_13), .dout_14(dout_5_14), .dout_15(dout_5_15), .dout_16(dout_5_16), .dout_17(dout_5_17), .dout_18(dout_5_18), .dout_19(dout_5_19), .dout_20(dout_5_20), .dout_21(dout_5_21), .dout_22(dout_5_22), .dout_23(dout_5_23), .dout_24(dout_5_24), .dout_25(dout_5_25), .dout_26(dout_5_26), .dout_27(dout_5_27), .dout_28(dout_5_28), .dout_29(dout_5_29), .dout_30(dout_5_30), .dout_31(dout_5_31), .dout_32(dout_5_32));
	SystolicBank # (.iWidth(iWidth), .oWidth(oWidth), .nRows(nRows), .nCols(nCols)) bank_6(.clk(clk), .rst(rst), .in_en(in_en), .config_load(pe_config_load), .iconfig_1(pe_config_6_1), .iconfig_2(pe_config_6_2), .iconfig_3(pe_config_6_3), .weight_1(weight_6_1), .weight_2(weight_6_2), .weight_3(weight_6_3), .feature_1(feature_1), .feature_2(feature_2), .feature_3(feature_3), .feature_4(feature_4), .feature_5(feature_5), .feature_6(feature_6), .feature_7(feature_7), .feature_8(feature_8), .feature_9(feature_9), .feature_10(feature_10), .feature_11(feature_11), .feature_12(feature_12), .feature_13(feature_13), .feature_14(feature_14), .feature_15(feature_15), .feature_16(feature_16), .feature_17(feature_17), .feature_18(feature_18), .feature_19(feature_19), .feature_20(feature_20), .feature_21(feature_21), .feature_22(feature_22), .feature_23(feature_23), .feature_24(feature_24), .feature_25(feature_25), .feature_26(feature_26), .feature_27(feature_27), .feature_28(feature_28), .feature_29(feature_29), .feature_30(feature_30), .feature_31(feature_31), .feature_32(feature_32), .feature_33(feature_33), .feature_34(feature_34), .A_1(A_1), .A_2(A_2), .A_3(A_3), .A_4(A_4), .A_5(A_5), .A_6(A_6), .A_7(A_7), .A_8(A_8), .A_9(A_9), .A_10(A_10), .A_11(A_11), .A_12(A_12), .A_13(A_13), .A_14(A_14), .A_15(A_15), .A_16(A_16), .A_17(A_17), .A_18(A_18), .A_19(A_19), .A_20(A_20), .A_21(A_21), .A_22(A_22), .A_23(A_23), .A_24(A_24), .A_25(A_25), .A_26(A_26), .A_27(A_27), .A_28(A_28), .A_29(A_29), .A_30(A_30), .A_31(A_31), .A_32(A_32), .B_1(B_1), .B_2(B_2), .B_3(B_3), .B_4(B_4), .B_5(B_5), .B_6(B_6), .B_7(B_7), .B_8(B_8), .B_9(B_9), .B_10(B_10), .B_11(B_11), .B_12(B_12), .B_13(B_13), .B_14(B_14), .B_15(B_15), .B_16(B_16), .B_17(B_17), .B_18(B_18), .B_19(B_19), .B_20(B_20), .B_21(B_21), .B_22(B_22), .B_23(B_23), .B_24(B_24), .B_25(B_25), .B_26(B_26), .B_27(B_27), .B_28(B_28), .B_29(B_29), .B_30(B_30), .B_31(B_31), .B_32(B_32), .C_1(C_1), .C_2(C_2), .C_3(C_3), .C_4(C_4), .C_5(C_5), .C_6(C_6), .C_7(C_7), .C_8(C_8), .C_9(C_9), .C_10(C_10), .C_11(C_11), .C_12(C_12), .C_13(C_13), .C_14(C_14), .C_15(C_15), .C_16(C_16), .C_17(C_17), .C_18(C_18), .C_19(C_19), .C_20(C_20), .C_21(C_21), .C_22(C_22), .C_23(C_23), .C_24(C_24), .C_25(C_25), .C_26(C_26), .C_27(C_27), .C_28(C_28), .C_29(C_29), .C_30(C_30), .C_31(C_31), .C_32(C_32), .D_1(D_1), .D_2(D_2), .D_3(D_3), .D_4(D_4), .D_5(D_5), .D_6(D_6), .D_7(D_7), .D_8(D_8), .D_9(D_9), .D_10(D_10), .D_11(D_11), .D_12(D_12), .D_13(D_13), .D_14(D_14), .D_15(D_15), .D_16(D_16), .D_17(D_17), .D_18(D_18), .D_19(D_19), .D_20(D_20), .D_21(D_21), .D_22(D_22), .D_23(D_23), .D_24(D_24), .D_25(D_25), .D_26(D_26), .D_27(D_27), .D_28(D_28), .D_29(D_29), .D_30(D_30), .D_31(D_31), .D_32(D_32), .E_1(E_1), .E_2(E_2), .E_3(E_3), .E_4(E_4), .E_5(E_5), .E_6(E_6), .E_7(E_7), .E_8(E_8), .E_9(E_9), .E_10(E_10), .E_11(E_11), .E_12(E_12), .E_13(E_13), .E_14(E_14), .E_15(E_15), .E_16(E_16), .E_17(E_17), .E_18(E_18), .E_19(E_19), .E_20(E_20), .E_21(E_21), .E_22(E_22), .E_23(E_23), .E_24(E_24), .E_25(E_25), .E_26(E_26), .E_27(E_27), .E_28(E_28), .E_29(E_29), .E_30(E_30), .E_31(E_31), .E_32(E_32), .F_1(F_1), .F_2(F_2), .F_3(F_3), .F_4(F_4), .F_5(F_5), .F_6(F_6), .F_7(F_7), .F_8(F_8), .F_9(F_9), .F_10(F_10), .F_11(F_11), .F_12(F_12), .F_13(F_13), .F_14(F_14), .F_15(F_15), .F_16(F_16), .F_17(F_17), .F_18(F_18), .F_19(F_19), .F_20(F_20), .F_21(F_21), .F_22(F_22), .F_23(F_23), .F_24(F_24), .F_25(F_25), .F_26(F_26), .F_27(F_27), .F_28(F_28), .F_29(F_29), .F_30(F_30), .F_31(F_31), .F_32(F_32), .G_1(G_1), .G_2(G_2), .G_3(G_3), .G_4(G_4), .G_5(G_5), .G_6(G_6), .G_7(G_7), .G_8(G_8), .G_9(G_9), .G_10(G_10), .G_11(G_11), .G_12(G_12), .G_13(G_13), .G_14(G_14), .G_15(G_15), .G_16(G_16), .G_17(G_17), .G_18(G_18), .G_19(G_19), .G_20(G_20), .G_21(G_21), .G_22(G_22), .G_23(G_23), .G_24(G_24), .G_25(G_25), .G_26(G_26), .G_27(G_27), .G_28(G_28), .G_29(G_29), .G_30(G_30), .G_31(G_31), .G_32(G_32), .dout_1(dout_6_1), .dout_2(dout_6_2), .dout_3(dout_6_3), .dout_4(dout_6_4), .dout_5(dout_6_5), .dout_6(dout_6_6), .dout_7(dout_6_7), .dout_8(dout_6_8), .dout_9(dout_6_9), .dout_10(dout_6_10), .dout_11(dout_6_11), .dout_12(dout_6_12), .dout_13(dout_6_13), .dout_14(dout_6_14), .dout_15(dout_6_15), .dout_16(dout_6_16), .dout_17(dout_6_17), .dout_18(dout_6_18), .dout_19(dout_6_19), .dout_20(dout_6_20), .dout_21(dout_6_21), .dout_22(dout_6_22), .dout_23(dout_6_23), .dout_24(dout_6_24), .dout_25(dout_6_25), .dout_26(dout_6_26), .dout_27(dout_6_27), .dout_28(dout_6_28), .dout_29(dout_6_29), .dout_30(dout_6_30), .dout_31(dout_6_31), .dout_32(dout_6_32));
	SystolicBank # (.iWidth(iWidth), .oWidth(oWidth), .nRows(nRows), .nCols(nCols)) bank_7(.clk(clk), .rst(rst), .in_en(in_en), .config_load(pe_config_load), .iconfig_1(pe_config_7_1), .iconfig_2(pe_config_7_2), .iconfig_3(pe_config_7_3), .weight_1(weight_7_1), .weight_2(weight_7_2), .weight_3(weight_7_3), .feature_1(feature_1), .feature_2(feature_2), .feature_3(feature_3), .feature_4(feature_4), .feature_5(feature_5), .feature_6(feature_6), .feature_7(feature_7), .feature_8(feature_8), .feature_9(feature_9), .feature_10(feature_10), .feature_11(feature_11), .feature_12(feature_12), .feature_13(feature_13), .feature_14(feature_14), .feature_15(feature_15), .feature_16(feature_16), .feature_17(feature_17), .feature_18(feature_18), .feature_19(feature_19), .feature_20(feature_20), .feature_21(feature_21), .feature_22(feature_22), .feature_23(feature_23), .feature_24(feature_24), .feature_25(feature_25), .feature_26(feature_26), .feature_27(feature_27), .feature_28(feature_28), .feature_29(feature_29), .feature_30(feature_30), .feature_31(feature_31), .feature_32(feature_32), .feature_33(feature_33), .feature_34(feature_34), .A_1(A_1), .A_2(A_2), .A_3(A_3), .A_4(A_4), .A_5(A_5), .A_6(A_6), .A_7(A_7), .A_8(A_8), .A_9(A_9), .A_10(A_10), .A_11(A_11), .A_12(A_12), .A_13(A_13), .A_14(A_14), .A_15(A_15), .A_16(A_16), .A_17(A_17), .A_18(A_18), .A_19(A_19), .A_20(A_20), .A_21(A_21), .A_22(A_22), .A_23(A_23), .A_24(A_24), .A_25(A_25), .A_26(A_26), .A_27(A_27), .A_28(A_28), .A_29(A_29), .A_30(A_30), .A_31(A_31), .A_32(A_32), .B_1(B_1), .B_2(B_2), .B_3(B_3), .B_4(B_4), .B_5(B_5), .B_6(B_6), .B_7(B_7), .B_8(B_8), .B_9(B_9), .B_10(B_10), .B_11(B_11), .B_12(B_12), .B_13(B_13), .B_14(B_14), .B_15(B_15), .B_16(B_16), .B_17(B_17), .B_18(B_18), .B_19(B_19), .B_20(B_20), .B_21(B_21), .B_22(B_22), .B_23(B_23), .B_24(B_24), .B_25(B_25), .B_26(B_26), .B_27(B_27), .B_28(B_28), .B_29(B_29), .B_30(B_30), .B_31(B_31), .B_32(B_32), .C_1(C_1), .C_2(C_2), .C_3(C_3), .C_4(C_4), .C_5(C_5), .C_6(C_6), .C_7(C_7), .C_8(C_8), .C_9(C_9), .C_10(C_10), .C_11(C_11), .C_12(C_12), .C_13(C_13), .C_14(C_14), .C_15(C_15), .C_16(C_16), .C_17(C_17), .C_18(C_18), .C_19(C_19), .C_20(C_20), .C_21(C_21), .C_22(C_22), .C_23(C_23), .C_24(C_24), .C_25(C_25), .C_26(C_26), .C_27(C_27), .C_28(C_28), .C_29(C_29), .C_30(C_30), .C_31(C_31), .C_32(C_32), .D_1(D_1), .D_2(D_2), .D_3(D_3), .D_4(D_4), .D_5(D_5), .D_6(D_6), .D_7(D_7), .D_8(D_8), .D_9(D_9), .D_10(D_10), .D_11(D_11), .D_12(D_12), .D_13(D_13), .D_14(D_14), .D_15(D_15), .D_16(D_16), .D_17(D_17), .D_18(D_18), .D_19(D_19), .D_20(D_20), .D_21(D_21), .D_22(D_22), .D_23(D_23), .D_24(D_24), .D_25(D_25), .D_26(D_26), .D_27(D_27), .D_28(D_28), .D_29(D_29), .D_30(D_30), .D_31(D_31), .D_32(D_32), .E_1(E_1), .E_2(E_2), .E_3(E_3), .E_4(E_4), .E_5(E_5), .E_6(E_6), .E_7(E_7), .E_8(E_8), .E_9(E_9), .E_10(E_10), .E_11(E_11), .E_12(E_12), .E_13(E_13), .E_14(E_14), .E_15(E_15), .E_16(E_16), .E_17(E_17), .E_18(E_18), .E_19(E_19), .E_20(E_20), .E_21(E_21), .E_22(E_22), .E_23(E_23), .E_24(E_24), .E_25(E_25), .E_26(E_26), .E_27(E_27), .E_28(E_28), .E_29(E_29), .E_30(E_30), .E_31(E_31), .E_32(E_32), .F_1(F_1), .F_2(F_2), .F_3(F_3), .F_4(F_4), .F_5(F_5), .F_6(F_6), .F_7(F_7), .F_8(F_8), .F_9(F_9), .F_10(F_10), .F_11(F_11), .F_12(F_12), .F_13(F_13), .F_14(F_14), .F_15(F_15), .F_16(F_16), .F_17(F_17), .F_18(F_18), .F_19(F_19), .F_20(F_20), .F_21(F_21), .F_22(F_22), .F_23(F_23), .F_24(F_24), .F_25(F_25), .F_26(F_26), .F_27(F_27), .F_28(F_28), .F_29(F_29), .F_30(F_30), .F_31(F_31), .F_32(F_32), .G_1(G_1), .G_2(G_2), .G_3(G_3), .G_4(G_4), .G_5(G_5), .G_6(G_6), .G_7(G_7), .G_8(G_8), .G_9(G_9), .G_10(G_10), .G_11(G_11), .G_12(G_12), .G_13(G_13), .G_14(G_14), .G_15(G_15), .G_16(G_16), .G_17(G_17), .G_18(G_18), .G_19(G_19), .G_20(G_20), .G_21(G_21), .G_22(G_22), .G_23(G_23), .G_24(G_24), .G_25(G_25), .G_26(G_26), .G_27(G_27), .G_28(G_28), .G_29(G_29), .G_30(G_30), .G_31(G_31), .G_32(G_32), .dout_1(dout_7_1), .dout_2(dout_7_2), .dout_3(dout_7_3), .dout_4(dout_7_4), .dout_5(dout_7_5), .dout_6(dout_7_6), .dout_7(dout_7_7), .dout_8(dout_7_8), .dout_9(dout_7_9), .dout_10(dout_7_10), .dout_11(dout_7_11), .dout_12(dout_7_12), .dout_13(dout_7_13), .dout_14(dout_7_14), .dout_15(dout_7_15), .dout_16(dout_7_16), .dout_17(dout_7_17), .dout_18(dout_7_18), .dout_19(dout_7_19), .dout_20(dout_7_20), .dout_21(dout_7_21), .dout_22(dout_7_22), .dout_23(dout_7_23), .dout_24(dout_7_24), .dout_25(dout_7_25), .dout_26(dout_7_26), .dout_27(dout_7_27), .dout_28(dout_7_28), .dout_29(dout_7_29), .dout_30(dout_7_30), .dout_31(dout_7_31), .dout_32(dout_7_32));
	SystolicBank # (.iWidth(iWidth), .oWidth(oWidth), .nRows(nRows), .nCols(nCols)) bank_8(.clk(clk), .rst(rst), .in_en(in_en), .config_load(pe_config_load), .iconfig_1(pe_config_8_1), .iconfig_2(pe_config_8_2), .iconfig_3(pe_config_8_3), .weight_1(weight_8_1), .weight_2(weight_8_2), .weight_3(weight_8_3), .feature_1(feature_1), .feature_2(feature_2), .feature_3(feature_3), .feature_4(feature_4), .feature_5(feature_5), .feature_6(feature_6), .feature_7(feature_7), .feature_8(feature_8), .feature_9(feature_9), .feature_10(feature_10), .feature_11(feature_11), .feature_12(feature_12), .feature_13(feature_13), .feature_14(feature_14), .feature_15(feature_15), .feature_16(feature_16), .feature_17(feature_17), .feature_18(feature_18), .feature_19(feature_19), .feature_20(feature_20), .feature_21(feature_21), .feature_22(feature_22), .feature_23(feature_23), .feature_24(feature_24), .feature_25(feature_25), .feature_26(feature_26), .feature_27(feature_27), .feature_28(feature_28), .feature_29(feature_29), .feature_30(feature_30), .feature_31(feature_31), .feature_32(feature_32), .feature_33(feature_33), .feature_34(feature_34), .A_1(A_1), .A_2(A_2), .A_3(A_3), .A_4(A_4), .A_5(A_5), .A_6(A_6), .A_7(A_7), .A_8(A_8), .A_9(A_9), .A_10(A_10), .A_11(A_11), .A_12(A_12), .A_13(A_13), .A_14(A_14), .A_15(A_15), .A_16(A_16), .A_17(A_17), .A_18(A_18), .A_19(A_19), .A_20(A_20), .A_21(A_21), .A_22(A_22), .A_23(A_23), .A_24(A_24), .A_25(A_25), .A_26(A_26), .A_27(A_27), .A_28(A_28), .A_29(A_29), .A_30(A_30), .A_31(A_31), .A_32(A_32), .B_1(B_1), .B_2(B_2), .B_3(B_3), .B_4(B_4), .B_5(B_5), .B_6(B_6), .B_7(B_7), .B_8(B_8), .B_9(B_9), .B_10(B_10), .B_11(B_11), .B_12(B_12), .B_13(B_13), .B_14(B_14), .B_15(B_15), .B_16(B_16), .B_17(B_17), .B_18(B_18), .B_19(B_19), .B_20(B_20), .B_21(B_21), .B_22(B_22), .B_23(B_23), .B_24(B_24), .B_25(B_25), .B_26(B_26), .B_27(B_27), .B_28(B_28), .B_29(B_29), .B_30(B_30), .B_31(B_31), .B_32(B_32), .C_1(C_1), .C_2(C_2), .C_3(C_3), .C_4(C_4), .C_5(C_5), .C_6(C_6), .C_7(C_7), .C_8(C_8), .C_9(C_9), .C_10(C_10), .C_11(C_11), .C_12(C_12), .C_13(C_13), .C_14(C_14), .C_15(C_15), .C_16(C_16), .C_17(C_17), .C_18(C_18), .C_19(C_19), .C_20(C_20), .C_21(C_21), .C_22(C_22), .C_23(C_23), .C_24(C_24), .C_25(C_25), .C_26(C_26), .C_27(C_27), .C_28(C_28), .C_29(C_29), .C_30(C_30), .C_31(C_31), .C_32(C_32), .D_1(D_1), .D_2(D_2), .D_3(D_3), .D_4(D_4), .D_5(D_5), .D_6(D_6), .D_7(D_7), .D_8(D_8), .D_9(D_9), .D_10(D_10), .D_11(D_11), .D_12(D_12), .D_13(D_13), .D_14(D_14), .D_15(D_15), .D_16(D_16), .D_17(D_17), .D_18(D_18), .D_19(D_19), .D_20(D_20), .D_21(D_21), .D_22(D_22), .D_23(D_23), .D_24(D_24), .D_25(D_25), .D_26(D_26), .D_27(D_27), .D_28(D_28), .D_29(D_29), .D_30(D_30), .D_31(D_31), .D_32(D_32), .E_1(E_1), .E_2(E_2), .E_3(E_3), .E_4(E_4), .E_5(E_5), .E_6(E_6), .E_7(E_7), .E_8(E_8), .E_9(E_9), .E_10(E_10), .E_11(E_11), .E_12(E_12), .E_13(E_13), .E_14(E_14), .E_15(E_15), .E_16(E_16), .E_17(E_17), .E_18(E_18), .E_19(E_19), .E_20(E_20), .E_21(E_21), .E_22(E_22), .E_23(E_23), .E_24(E_24), .E_25(E_25), .E_26(E_26), .E_27(E_27), .E_28(E_28), .E_29(E_29), .E_30(E_30), .E_31(E_31), .E_32(E_32), .F_1(F_1), .F_2(F_2), .F_3(F_3), .F_4(F_4), .F_5(F_5), .F_6(F_6), .F_7(F_7), .F_8(F_8), .F_9(F_9), .F_10(F_10), .F_11(F_11), .F_12(F_12), .F_13(F_13), .F_14(F_14), .F_15(F_15), .F_16(F_16), .F_17(F_17), .F_18(F_18), .F_19(F_19), .F_20(F_20), .F_21(F_21), .F_22(F_22), .F_23(F_23), .F_24(F_24), .F_25(F_25), .F_26(F_26), .F_27(F_27), .F_28(F_28), .F_29(F_29), .F_30(F_30), .F_31(F_31), .F_32(F_32), .G_1(G_1), .G_2(G_2), .G_3(G_3), .G_4(G_4), .G_5(G_5), .G_6(G_6), .G_7(G_7), .G_8(G_8), .G_9(G_9), .G_10(G_10), .G_11(G_11), .G_12(G_12), .G_13(G_13), .G_14(G_14), .G_15(G_15), .G_16(G_16), .G_17(G_17), .G_18(G_18), .G_19(G_19), .G_20(G_20), .G_21(G_21), .G_22(G_22), .G_23(G_23), .G_24(G_24), .G_25(G_25), .G_26(G_26), .G_27(G_27), .G_28(G_28), .G_29(G_29), .G_30(G_30), .G_31(G_31), .G_32(G_32), .dout_1(dout_8_1), .dout_2(dout_8_2), .dout_3(dout_8_3), .dout_4(dout_8_4), .dout_5(dout_8_5), .dout_6(dout_8_6), .dout_7(dout_8_7), .dout_8(dout_8_8), .dout_9(dout_8_9), .dout_10(dout_8_10), .dout_11(dout_8_11), .dout_12(dout_8_12), .dout_13(dout_8_13), .dout_14(dout_8_14), .dout_15(dout_8_15), .dout_16(dout_8_16), .dout_17(dout_8_17), .dout_18(dout_8_18), .dout_19(dout_8_19), .dout_20(dout_8_20), .dout_21(dout_8_21), .dout_22(dout_8_22), .dout_23(dout_8_23), .dout_24(dout_8_24), .dout_25(dout_8_25), .dout_26(dout_8_26), .dout_27(dout_8_27), .dout_28(dout_8_28), .dout_29(dout_8_29), .dout_30(dout_8_30), .dout_31(dout_8_31), .dout_32(dout_8_32));
	SystolicBank # (.iWidth(iWidth), .oWidth(oWidth), .nRows(nRows), .nCols(nCols)) bank_9(.clk(clk), .rst(rst), .in_en(in_en), .config_load(pe_config_load), .iconfig_1(pe_config_9_1), .iconfig_2(pe_config_9_2), .iconfig_3(pe_config_9_3), .weight_1(weight_9_1), .weight_2(weight_9_2), .weight_3(weight_9_3), .feature_1(feature_1), .feature_2(feature_2), .feature_3(feature_3), .feature_4(feature_4), .feature_5(feature_5), .feature_6(feature_6), .feature_7(feature_7), .feature_8(feature_8), .feature_9(feature_9), .feature_10(feature_10), .feature_11(feature_11), .feature_12(feature_12), .feature_13(feature_13), .feature_14(feature_14), .feature_15(feature_15), .feature_16(feature_16), .feature_17(feature_17), .feature_18(feature_18), .feature_19(feature_19), .feature_20(feature_20), .feature_21(feature_21), .feature_22(feature_22), .feature_23(feature_23), .feature_24(feature_24), .feature_25(feature_25), .feature_26(feature_26), .feature_27(feature_27), .feature_28(feature_28), .feature_29(feature_29), .feature_30(feature_30), .feature_31(feature_31), .feature_32(feature_32), .feature_33(feature_33), .feature_34(feature_34), .A_1(A_1), .A_2(A_2), .A_3(A_3), .A_4(A_4), .A_5(A_5), .A_6(A_6), .A_7(A_7), .A_8(A_8), .A_9(A_9), .A_10(A_10), .A_11(A_11), .A_12(A_12), .A_13(A_13), .A_14(A_14), .A_15(A_15), .A_16(A_16), .A_17(A_17), .A_18(A_18), .A_19(A_19), .A_20(A_20), .A_21(A_21), .A_22(A_22), .A_23(A_23), .A_24(A_24), .A_25(A_25), .A_26(A_26), .A_27(A_27), .A_28(A_28), .A_29(A_29), .A_30(A_30), .A_31(A_31), .A_32(A_32), .B_1(B_1), .B_2(B_2), .B_3(B_3), .B_4(B_4), .B_5(B_5), .B_6(B_6), .B_7(B_7), .B_8(B_8), .B_9(B_9), .B_10(B_10), .B_11(B_11), .B_12(B_12), .B_13(B_13), .B_14(B_14), .B_15(B_15), .B_16(B_16), .B_17(B_17), .B_18(B_18), .B_19(B_19), .B_20(B_20), .B_21(B_21), .B_22(B_22), .B_23(B_23), .B_24(B_24), .B_25(B_25), .B_26(B_26), .B_27(B_27), .B_28(B_28), .B_29(B_29), .B_30(B_30), .B_31(B_31), .B_32(B_32), .C_1(C_1), .C_2(C_2), .C_3(C_3), .C_4(C_4), .C_5(C_5), .C_6(C_6), .C_7(C_7), .C_8(C_8), .C_9(C_9), .C_10(C_10), .C_11(C_11), .C_12(C_12), .C_13(C_13), .C_14(C_14), .C_15(C_15), .C_16(C_16), .C_17(C_17), .C_18(C_18), .C_19(C_19), .C_20(C_20), .C_21(C_21), .C_22(C_22), .C_23(C_23), .C_24(C_24), .C_25(C_25), .C_26(C_26), .C_27(C_27), .C_28(C_28), .C_29(C_29), .C_30(C_30), .C_31(C_31), .C_32(C_32), .D_1(D_1), .D_2(D_2), .D_3(D_3), .D_4(D_4), .D_5(D_5), .D_6(D_6), .D_7(D_7), .D_8(D_8), .D_9(D_9), .D_10(D_10), .D_11(D_11), .D_12(D_12), .D_13(D_13), .D_14(D_14), .D_15(D_15), .D_16(D_16), .D_17(D_17), .D_18(D_18), .D_19(D_19), .D_20(D_20), .D_21(D_21), .D_22(D_22), .D_23(D_23), .D_24(D_24), .D_25(D_25), .D_26(D_26), .D_27(D_27), .D_28(D_28), .D_29(D_29), .D_30(D_30), .D_31(D_31), .D_32(D_32), .E_1(E_1), .E_2(E_2), .E_3(E_3), .E_4(E_4), .E_5(E_5), .E_6(E_6), .E_7(E_7), .E_8(E_8), .E_9(E_9), .E_10(E_10), .E_11(E_11), .E_12(E_12), .E_13(E_13), .E_14(E_14), .E_15(E_15), .E_16(E_16), .E_17(E_17), .E_18(E_18), .E_19(E_19), .E_20(E_20), .E_21(E_21), .E_22(E_22), .E_23(E_23), .E_24(E_24), .E_25(E_25), .E_26(E_26), .E_27(E_27), .E_28(E_28), .E_29(E_29), .E_30(E_30), .E_31(E_31), .E_32(E_32), .F_1(F_1), .F_2(F_2), .F_3(F_3), .F_4(F_4), .F_5(F_5), .F_6(F_6), .F_7(F_7), .F_8(F_8), .F_9(F_9), .F_10(F_10), .F_11(F_11), .F_12(F_12), .F_13(F_13), .F_14(F_14), .F_15(F_15), .F_16(F_16), .F_17(F_17), .F_18(F_18), .F_19(F_19), .F_20(F_20), .F_21(F_21), .F_22(F_22), .F_23(F_23), .F_24(F_24), .F_25(F_25), .F_26(F_26), .F_27(F_27), .F_28(F_28), .F_29(F_29), .F_30(F_30), .F_31(F_31), .F_32(F_32), .G_1(G_1), .G_2(G_2), .G_3(G_3), .G_4(G_4), .G_5(G_5), .G_6(G_6), .G_7(G_7), .G_8(G_8), .G_9(G_9), .G_10(G_10), .G_11(G_11), .G_12(G_12), .G_13(G_13), .G_14(G_14), .G_15(G_15), .G_16(G_16), .G_17(G_17), .G_18(G_18), .G_19(G_19), .G_20(G_20), .G_21(G_21), .G_22(G_22), .G_23(G_23), .G_24(G_24), .G_25(G_25), .G_26(G_26), .G_27(G_27), .G_28(G_28), .G_29(G_29), .G_30(G_30), .G_31(G_31), .G_32(G_32), .dout_1(dout_9_1), .dout_2(dout_9_2), .dout_3(dout_9_3), .dout_4(dout_9_4), .dout_5(dout_9_5), .dout_6(dout_9_6), .dout_7(dout_9_7), .dout_8(dout_9_8), .dout_9(dout_9_9), .dout_10(dout_9_10), .dout_11(dout_9_11), .dout_12(dout_9_12), .dout_13(dout_9_13), .dout_14(dout_9_14), .dout_15(dout_9_15), .dout_16(dout_9_16), .dout_17(dout_9_17), .dout_18(dout_9_18), .dout_19(dout_9_19), .dout_20(dout_9_20), .dout_21(dout_9_21), .dout_22(dout_9_22), .dout_23(dout_9_23), .dout_24(dout_9_24), .dout_25(dout_9_25), .dout_26(dout_9_26), .dout_27(dout_9_27), .dout_28(dout_9_28), .dout_29(dout_9_29), .dout_30(dout_9_30), .dout_31(dout_9_31), .dout_32(dout_9_32));
	SystolicBank # (.iWidth(iWidth), .oWidth(oWidth), .nRows(nRows), .nCols(nCols)) bank_10(.clk(clk), .rst(rst), .in_en(in_en), .config_load(pe_config_load), .iconfig_1(pe_config_10_1), .iconfig_2(pe_config_10_2), .iconfig_3(pe_config_10_3), .weight_1(weight_10_1), .weight_2(weight_10_2), .weight_3(weight_10_3), .feature_1(feature_1), .feature_2(feature_2), .feature_3(feature_3), .feature_4(feature_4), .feature_5(feature_5), .feature_6(feature_6), .feature_7(feature_7), .feature_8(feature_8), .feature_9(feature_9), .feature_10(feature_10), .feature_11(feature_11), .feature_12(feature_12), .feature_13(feature_13), .feature_14(feature_14), .feature_15(feature_15), .feature_16(feature_16), .feature_17(feature_17), .feature_18(feature_18), .feature_19(feature_19), .feature_20(feature_20), .feature_21(feature_21), .feature_22(feature_22), .feature_23(feature_23), .feature_24(feature_24), .feature_25(feature_25), .feature_26(feature_26), .feature_27(feature_27), .feature_28(feature_28), .feature_29(feature_29), .feature_30(feature_30), .feature_31(feature_31), .feature_32(feature_32), .feature_33(feature_33), .feature_34(feature_34), .A_1(A_1), .A_2(A_2), .A_3(A_3), .A_4(A_4), .A_5(A_5), .A_6(A_6), .A_7(A_7), .A_8(A_8), .A_9(A_9), .A_10(A_10), .A_11(A_11), .A_12(A_12), .A_13(A_13), .A_14(A_14), .A_15(A_15), .A_16(A_16), .A_17(A_17), .A_18(A_18), .A_19(A_19), .A_20(A_20), .A_21(A_21), .A_22(A_22), .A_23(A_23), .A_24(A_24), .A_25(A_25), .A_26(A_26), .A_27(A_27), .A_28(A_28), .A_29(A_29), .A_30(A_30), .A_31(A_31), .A_32(A_32), .B_1(B_1), .B_2(B_2), .B_3(B_3), .B_4(B_4), .B_5(B_5), .B_6(B_6), .B_7(B_7), .B_8(B_8), .B_9(B_9), .B_10(B_10), .B_11(B_11), .B_12(B_12), .B_13(B_13), .B_14(B_14), .B_15(B_15), .B_16(B_16), .B_17(B_17), .B_18(B_18), .B_19(B_19), .B_20(B_20), .B_21(B_21), .B_22(B_22), .B_23(B_23), .B_24(B_24), .B_25(B_25), .B_26(B_26), .B_27(B_27), .B_28(B_28), .B_29(B_29), .B_30(B_30), .B_31(B_31), .B_32(B_32), .C_1(C_1), .C_2(C_2), .C_3(C_3), .C_4(C_4), .C_5(C_5), .C_6(C_6), .C_7(C_7), .C_8(C_8), .C_9(C_9), .C_10(C_10), .C_11(C_11), .C_12(C_12), .C_13(C_13), .C_14(C_14), .C_15(C_15), .C_16(C_16), .C_17(C_17), .C_18(C_18), .C_19(C_19), .C_20(C_20), .C_21(C_21), .C_22(C_22), .C_23(C_23), .C_24(C_24), .C_25(C_25), .C_26(C_26), .C_27(C_27), .C_28(C_28), .C_29(C_29), .C_30(C_30), .C_31(C_31), .C_32(C_32), .D_1(D_1), .D_2(D_2), .D_3(D_3), .D_4(D_4), .D_5(D_5), .D_6(D_6), .D_7(D_7), .D_8(D_8), .D_9(D_9), .D_10(D_10), .D_11(D_11), .D_12(D_12), .D_13(D_13), .D_14(D_14), .D_15(D_15), .D_16(D_16), .D_17(D_17), .D_18(D_18), .D_19(D_19), .D_20(D_20), .D_21(D_21), .D_22(D_22), .D_23(D_23), .D_24(D_24), .D_25(D_25), .D_26(D_26), .D_27(D_27), .D_28(D_28), .D_29(D_29), .D_30(D_30), .D_31(D_31), .D_32(D_32), .E_1(E_1), .E_2(E_2), .E_3(E_3), .E_4(E_4), .E_5(E_5), .E_6(E_6), .E_7(E_7), .E_8(E_8), .E_9(E_9), .E_10(E_10), .E_11(E_11), .E_12(E_12), .E_13(E_13), .E_14(E_14), .E_15(E_15), .E_16(E_16), .E_17(E_17), .E_18(E_18), .E_19(E_19), .E_20(E_20), .E_21(E_21), .E_22(E_22), .E_23(E_23), .E_24(E_24), .E_25(E_25), .E_26(E_26), .E_27(E_27), .E_28(E_28), .E_29(E_29), .E_30(E_30), .E_31(E_31), .E_32(E_32), .F_1(F_1), .F_2(F_2), .F_3(F_3), .F_4(F_4), .F_5(F_5), .F_6(F_6), .F_7(F_7), .F_8(F_8), .F_9(F_9), .F_10(F_10), .F_11(F_11), .F_12(F_12), .F_13(F_13), .F_14(F_14), .F_15(F_15), .F_16(F_16), .F_17(F_17), .F_18(F_18), .F_19(F_19), .F_20(F_20), .F_21(F_21), .F_22(F_22), .F_23(F_23), .F_24(F_24), .F_25(F_25), .F_26(F_26), .F_27(F_27), .F_28(F_28), .F_29(F_29), .F_30(F_30), .F_31(F_31), .F_32(F_32), .G_1(G_1), .G_2(G_2), .G_3(G_3), .G_4(G_4), .G_5(G_5), .G_6(G_6), .G_7(G_7), .G_8(G_8), .G_9(G_9), .G_10(G_10), .G_11(G_11), .G_12(G_12), .G_13(G_13), .G_14(G_14), .G_15(G_15), .G_16(G_16), .G_17(G_17), .G_18(G_18), .G_19(G_19), .G_20(G_20), .G_21(G_21), .G_22(G_22), .G_23(G_23), .G_24(G_24), .G_25(G_25), .G_26(G_26), .G_27(G_27), .G_28(G_28), .G_29(G_29), .G_30(G_30), .G_31(G_31), .G_32(G_32), .dout_1(dout_10_1), .dout_2(dout_10_2), .dout_3(dout_10_3), .dout_4(dout_10_4), .dout_5(dout_10_5), .dout_6(dout_10_6), .dout_7(dout_10_7), .dout_8(dout_10_8), .dout_9(dout_10_9), .dout_10(dout_10_10), .dout_11(dout_10_11), .dout_12(dout_10_12), .dout_13(dout_10_13), .dout_14(dout_10_14), .dout_15(dout_10_15), .dout_16(dout_10_16), .dout_17(dout_10_17), .dout_18(dout_10_18), .dout_19(dout_10_19), .dout_20(dout_10_20), .dout_21(dout_10_21), .dout_22(dout_10_22), .dout_23(dout_10_23), .dout_24(dout_10_24), .dout_25(dout_10_25), .dout_26(dout_10_26), .dout_27(dout_10_27), .dout_28(dout_10_28), .dout_29(dout_10_29), .dout_30(dout_10_30), .dout_31(dout_10_31), .dout_32(dout_10_32));
	SystolicBank # (.iWidth(iWidth), .oWidth(oWidth), .nRows(nRows), .nCols(nCols)) bank_11(.clk(clk), .rst(rst), .in_en(in_en), .config_load(pe_config_load), .iconfig_1(pe_config_11_1), .iconfig_2(pe_config_11_2), .iconfig_3(pe_config_11_3), .weight_1(weight_11_1), .weight_2(weight_11_2), .weight_3(weight_11_3), .feature_1(feature_1), .feature_2(feature_2), .feature_3(feature_3), .feature_4(feature_4), .feature_5(feature_5), .feature_6(feature_6), .feature_7(feature_7), .feature_8(feature_8), .feature_9(feature_9), .feature_10(feature_10), .feature_11(feature_11), .feature_12(feature_12), .feature_13(feature_13), .feature_14(feature_14), .feature_15(feature_15), .feature_16(feature_16), .feature_17(feature_17), .feature_18(feature_18), .feature_19(feature_19), .feature_20(feature_20), .feature_21(feature_21), .feature_22(feature_22), .feature_23(feature_23), .feature_24(feature_24), .feature_25(feature_25), .feature_26(feature_26), .feature_27(feature_27), .feature_28(feature_28), .feature_29(feature_29), .feature_30(feature_30), .feature_31(feature_31), .feature_32(feature_32), .feature_33(feature_33), .feature_34(feature_34), .A_1(A_1), .A_2(A_2), .A_3(A_3), .A_4(A_4), .A_5(A_5), .A_6(A_6), .A_7(A_7), .A_8(A_8), .A_9(A_9), .A_10(A_10), .A_11(A_11), .A_12(A_12), .A_13(A_13), .A_14(A_14), .A_15(A_15), .A_16(A_16), .A_17(A_17), .A_18(A_18), .A_19(A_19), .A_20(A_20), .A_21(A_21), .A_22(A_22), .A_23(A_23), .A_24(A_24), .A_25(A_25), .A_26(A_26), .A_27(A_27), .A_28(A_28), .A_29(A_29), .A_30(A_30), .A_31(A_31), .A_32(A_32), .B_1(B_1), .B_2(B_2), .B_3(B_3), .B_4(B_4), .B_5(B_5), .B_6(B_6), .B_7(B_7), .B_8(B_8), .B_9(B_9), .B_10(B_10), .B_11(B_11), .B_12(B_12), .B_13(B_13), .B_14(B_14), .B_15(B_15), .B_16(B_16), .B_17(B_17), .B_18(B_18), .B_19(B_19), .B_20(B_20), .B_21(B_21), .B_22(B_22), .B_23(B_23), .B_24(B_24), .B_25(B_25), .B_26(B_26), .B_27(B_27), .B_28(B_28), .B_29(B_29), .B_30(B_30), .B_31(B_31), .B_32(B_32), .C_1(C_1), .C_2(C_2), .C_3(C_3), .C_4(C_4), .C_5(C_5), .C_6(C_6), .C_7(C_7), .C_8(C_8), .C_9(C_9), .C_10(C_10), .C_11(C_11), .C_12(C_12), .C_13(C_13), .C_14(C_14), .C_15(C_15), .C_16(C_16), .C_17(C_17), .C_18(C_18), .C_19(C_19), .C_20(C_20), .C_21(C_21), .C_22(C_22), .C_23(C_23), .C_24(C_24), .C_25(C_25), .C_26(C_26), .C_27(C_27), .C_28(C_28), .C_29(C_29), .C_30(C_30), .C_31(C_31), .C_32(C_32), .D_1(D_1), .D_2(D_2), .D_3(D_3), .D_4(D_4), .D_5(D_5), .D_6(D_6), .D_7(D_7), .D_8(D_8), .D_9(D_9), .D_10(D_10), .D_11(D_11), .D_12(D_12), .D_13(D_13), .D_14(D_14), .D_15(D_15), .D_16(D_16), .D_17(D_17), .D_18(D_18), .D_19(D_19), .D_20(D_20), .D_21(D_21), .D_22(D_22), .D_23(D_23), .D_24(D_24), .D_25(D_25), .D_26(D_26), .D_27(D_27), .D_28(D_28), .D_29(D_29), .D_30(D_30), .D_31(D_31), .D_32(D_32), .E_1(E_1), .E_2(E_2), .E_3(E_3), .E_4(E_4), .E_5(E_5), .E_6(E_6), .E_7(E_7), .E_8(E_8), .E_9(E_9), .E_10(E_10), .E_11(E_11), .E_12(E_12), .E_13(E_13), .E_14(E_14), .E_15(E_15), .E_16(E_16), .E_17(E_17), .E_18(E_18), .E_19(E_19), .E_20(E_20), .E_21(E_21), .E_22(E_22), .E_23(E_23), .E_24(E_24), .E_25(E_25), .E_26(E_26), .E_27(E_27), .E_28(E_28), .E_29(E_29), .E_30(E_30), .E_31(E_31), .E_32(E_32), .F_1(F_1), .F_2(F_2), .F_3(F_3), .F_4(F_4), .F_5(F_5), .F_6(F_6), .F_7(F_7), .F_8(F_8), .F_9(F_9), .F_10(F_10), .F_11(F_11), .F_12(F_12), .F_13(F_13), .F_14(F_14), .F_15(F_15), .F_16(F_16), .F_17(F_17), .F_18(F_18), .F_19(F_19), .F_20(F_20), .F_21(F_21), .F_22(F_22), .F_23(F_23), .F_24(F_24), .F_25(F_25), .F_26(F_26), .F_27(F_27), .F_28(F_28), .F_29(F_29), .F_30(F_30), .F_31(F_31), .F_32(F_32), .G_1(G_1), .G_2(G_2), .G_3(G_3), .G_4(G_4), .G_5(G_5), .G_6(G_6), .G_7(G_7), .G_8(G_8), .G_9(G_9), .G_10(G_10), .G_11(G_11), .G_12(G_12), .G_13(G_13), .G_14(G_14), .G_15(G_15), .G_16(G_16), .G_17(G_17), .G_18(G_18), .G_19(G_19), .G_20(G_20), .G_21(G_21), .G_22(G_22), .G_23(G_23), .G_24(G_24), .G_25(G_25), .G_26(G_26), .G_27(G_27), .G_28(G_28), .G_29(G_29), .G_30(G_30), .G_31(G_31), .G_32(G_32), .dout_1(dout_11_1), .dout_2(dout_11_2), .dout_3(dout_11_3), .dout_4(dout_11_4), .dout_5(dout_11_5), .dout_6(dout_11_6), .dout_7(dout_11_7), .dout_8(dout_11_8), .dout_9(dout_11_9), .dout_10(dout_11_10), .dout_11(dout_11_11), .dout_12(dout_11_12), .dout_13(dout_11_13), .dout_14(dout_11_14), .dout_15(dout_11_15), .dout_16(dout_11_16), .dout_17(dout_11_17), .dout_18(dout_11_18), .dout_19(dout_11_19), .dout_20(dout_11_20), .dout_21(dout_11_21), .dout_22(dout_11_22), .dout_23(dout_11_23), .dout_24(dout_11_24), .dout_25(dout_11_25), .dout_26(dout_11_26), .dout_27(dout_11_27), .dout_28(dout_11_28), .dout_29(dout_11_29), .dout_30(dout_11_30), .dout_31(dout_11_31), .dout_32(dout_11_32));

	DFSM # (.MAX_nPERIOD(MAX_nPERIOD), .MAX_nLMAC(MAX_nLMAC), .MAX_nSHFT(MAX_nSHFT)) fsm_1(.clk(clk), .rst(rst), .config_en(dfsm_config_en), .iconfig(dfsm_config), .in_en(in_en), .start(start), .in_en_bypass(dfsm_data_en_1), .out_en(dout_en_1), .start_out(start_bypass_1), .A(A_1), .B(B_1), .C(C_1), .D(D_1), .E(E_1), .F(F_1), .G(G_1));
	DFSM # (.MAX_nPERIOD(MAX_nPERIOD), .MAX_nLMAC(MAX_nLMAC), .MAX_nSHFT(MAX_nSHFT)) fsm_2(.clk(clk), .rst(rst), .config_en(dfsm_config_en), .iconfig(dfsm_config), .in_en(dfsm_data_en_1), .start(start_bypass_1), .in_en_bypass(dfsm_data_en_2), .out_en(dout_en_2), .start_out(start_bypass_2), .A(A_2), .B(B_2), .C(C_2), .D(D_2), .E(E_2), .F(F_2), .G(G_2));
	DFSM # (.MAX_nPERIOD(MAX_nPERIOD), .MAX_nLMAC(MAX_nLMAC), .MAX_nSHFT(MAX_nSHFT)) fsm_3(.clk(clk), .rst(rst), .config_en(dfsm_config_en), .iconfig(dfsm_config), .in_en(dfsm_data_en_2), .start(start_bypass_2), .in_en_bypass(dfsm_data_en_3), .out_en(dout_en_3), .start_out(start_bypass_3), .A(A_3), .B(B_3), .C(C_3), .D(D_3), .E(E_3), .F(F_3), .G(G_3));
	DFSM # (.MAX_nPERIOD(MAX_nPERIOD), .MAX_nLMAC(MAX_nLMAC), .MAX_nSHFT(MAX_nSHFT)) fsm_4(.clk(clk), .rst(rst), .config_en(dfsm_config_en), .iconfig(dfsm_config), .in_en(dfsm_data_en_3), .start(start_bypass_3), .in_en_bypass(dfsm_data_en_4), .out_en(dout_en_4), .start_out(start_bypass_4), .A(A_4), .B(B_4), .C(C_4), .D(D_4), .E(E_4), .F(F_4), .G(G_4));
	DFSM # (.MAX_nPERIOD(MAX_nPERIOD), .MAX_nLMAC(MAX_nLMAC), .MAX_nSHFT(MAX_nSHFT)) fsm_5(.clk(clk), .rst(rst), .config_en(dfsm_config_en), .iconfig(dfsm_config), .in_en(dfsm_data_en_4), .start(start_bypass_4), .in_en_bypass(dfsm_data_en_5), .out_en(dout_en_5), .start_out(start_bypass_5), .A(A_5), .B(B_5), .C(C_5), .D(D_5), .E(E_5), .F(F_5), .G(G_5));
	DFSM # (.MAX_nPERIOD(MAX_nPERIOD), .MAX_nLMAC(MAX_nLMAC), .MAX_nSHFT(MAX_nSHFT)) fsm_6(.clk(clk), .rst(rst), .config_en(dfsm_config_en), .iconfig(dfsm_config), .in_en(dfsm_data_en_5), .start(start_bypass_5), .in_en_bypass(dfsm_data_en_6), .out_en(dout_en_6), .start_out(start_bypass_6), .A(A_6), .B(B_6), .C(C_6), .D(D_6), .E(E_6), .F(F_6), .G(G_6));
	DFSM # (.MAX_nPERIOD(MAX_nPERIOD), .MAX_nLMAC(MAX_nLMAC), .MAX_nSHFT(MAX_nSHFT)) fsm_7(.clk(clk), .rst(rst), .config_en(dfsm_config_en), .iconfig(dfsm_config), .in_en(dfsm_data_en_6), .start(start_bypass_6), .in_en_bypass(dfsm_data_en_7), .out_en(dout_en_7), .start_out(start_bypass_7), .A(A_7), .B(B_7), .C(C_7), .D(D_7), .E(E_7), .F(F_7), .G(G_7));
	DFSM # (.MAX_nPERIOD(MAX_nPERIOD), .MAX_nLMAC(MAX_nLMAC), .MAX_nSHFT(MAX_nSHFT)) fsm_8(.clk(clk), .rst(rst), .config_en(dfsm_config_en), .iconfig(dfsm_config), .in_en(dfsm_data_en_7), .start(start_bypass_7), .in_en_bypass(dfsm_data_en_8), .out_en(dout_en_8), .start_out(start_bypass_8), .A(A_8), .B(B_8), .C(C_8), .D(D_8), .E(E_8), .F(F_8), .G(G_8));
	DFSM # (.MAX_nPERIOD(MAX_nPERIOD), .MAX_nLMAC(MAX_nLMAC), .MAX_nSHFT(MAX_nSHFT)) fsm_9(.clk(clk), .rst(rst), .config_en(dfsm_config_en), .iconfig(dfsm_config), .in_en(dfsm_data_en_8), .start(start_bypass_8), .in_en_bypass(dfsm_data_en_9), .out_en(dout_en_9), .start_out(start_bypass_9), .A(A_9), .B(B_9), .C(C_9), .D(D_9), .E(E_9), .F(F_9), .G(G_9));
	DFSM # (.MAX_nPERIOD(MAX_nPERIOD), .MAX_nLMAC(MAX_nLMAC), .MAX_nSHFT(MAX_nSHFT)) fsm_10(.clk(clk), .rst(rst), .config_en(dfsm_config_en), .iconfig(dfsm_config), .in_en(dfsm_data_en_9), .start(start_bypass_9), .in_en_bypass(dfsm_data_en_10), .out_en(dout_en_10), .start_out(start_bypass_10), .A(A_10), .B(B_10), .C(C_10), .D(D_10), .E(E_10), .F(F_10), .G(G_10));
	DFSM # (.MAX_nPERIOD(MAX_nPERIOD), .MAX_nLMAC(MAX_nLMAC), .MAX_nSHFT(MAX_nSHFT)) fsm_11(.clk(clk), .rst(rst), .config_en(dfsm_config_en), .iconfig(dfsm_config), .in_en(dfsm_data_en_10), .start(start_bypass_10), .in_en_bypass(dfsm_data_en_11), .out_en(dout_en_11), .start_out(start_bypass_11), .A(A_11), .B(B_11), .C(C_11), .D(D_11), .E(E_11), .F(F_11), .G(G_11));
	DFSM # (.MAX_nPERIOD(MAX_nPERIOD), .MAX_nLMAC(MAX_nLMAC), .MAX_nSHFT(MAX_nSHFT)) fsm_12(.clk(clk), .rst(rst), .config_en(dfsm_config_en), .iconfig(dfsm_config), .in_en(dfsm_data_en_11), .start(start_bypass_11), .in_en_bypass(dfsm_data_en_12), .out_en(dout_en_12), .start_out(start_bypass_12), .A(A_12), .B(B_12), .C(C_12), .D(D_12), .E(E_12), .F(F_12), .G(G_12));
	DFSM # (.MAX_nPERIOD(MAX_nPERIOD), .MAX_nLMAC(MAX_nLMAC), .MAX_nSHFT(MAX_nSHFT)) fsm_13(.clk(clk), .rst(rst), .config_en(dfsm_config_en), .iconfig(dfsm_config), .in_en(dfsm_data_en_12), .start(start_bypass_12), .in_en_bypass(dfsm_data_en_13), .out_en(dout_en_13), .start_out(start_bypass_13), .A(A_13), .B(B_13), .C(C_13), .D(D_13), .E(E_13), .F(F_13), .G(G_13));
	DFSM # (.MAX_nPERIOD(MAX_nPERIOD), .MAX_nLMAC(MAX_nLMAC), .MAX_nSHFT(MAX_nSHFT)) fsm_14(.clk(clk), .rst(rst), .config_en(dfsm_config_en), .iconfig(dfsm_config), .in_en(dfsm_data_en_13), .start(start_bypass_13), .in_en_bypass(dfsm_data_en_14), .out_en(dout_en_14), .start_out(start_bypass_14), .A(A_14), .B(B_14), .C(C_14), .D(D_14), .E(E_14), .F(F_14), .G(G_14));
	DFSM # (.MAX_nPERIOD(MAX_nPERIOD), .MAX_nLMAC(MAX_nLMAC), .MAX_nSHFT(MAX_nSHFT)) fsm_15(.clk(clk), .rst(rst), .config_en(dfsm_config_en), .iconfig(dfsm_config), .in_en(dfsm_data_en_14), .start(start_bypass_14), .in_en_bypass(dfsm_data_en_15), .out_en(dout_en_15), .start_out(start_bypass_15), .A(A_15), .B(B_15), .C(C_15), .D(D_15), .E(E_15), .F(F_15), .G(G_15));
	DFSM # (.MAX_nPERIOD(MAX_nPERIOD), .MAX_nLMAC(MAX_nLMAC), .MAX_nSHFT(MAX_nSHFT)) fsm_16(.clk(clk), .rst(rst), .config_en(dfsm_config_en), .iconfig(dfsm_config), .in_en(dfsm_data_en_15), .start(start_bypass_15), .in_en_bypass(dfsm_data_en_16), .out_en(dout_en_16), .start_out(start_bypass_16), .A(A_16), .B(B_16), .C(C_16), .D(D_16), .E(E_16), .F(F_16), .G(G_16));
	DFSM # (.MAX_nPERIOD(MAX_nPERIOD), .MAX_nLMAC(MAX_nLMAC), .MAX_nSHFT(MAX_nSHFT)) fsm_17(.clk(clk), .rst(rst), .config_en(dfsm_config_en), .iconfig(dfsm_config), .in_en(dfsm_data_en_16), .start(start_bypass_16), .in_en_bypass(dfsm_data_en_17), .out_en(dout_en_17), .start_out(start_bypass_17), .A(A_17), .B(B_17), .C(C_17), .D(D_17), .E(E_17), .F(F_17), .G(G_17));
	DFSM # (.MAX_nPERIOD(MAX_nPERIOD), .MAX_nLMAC(MAX_nLMAC), .MAX_nSHFT(MAX_nSHFT)) fsm_18(.clk(clk), .rst(rst), .config_en(dfsm_config_en), .iconfig(dfsm_config), .in_en(dfsm_data_en_17), .start(start_bypass_17), .in_en_bypass(dfsm_data_en_18), .out_en(dout_en_18), .start_out(start_bypass_18), .A(A_18), .B(B_18), .C(C_18), .D(D_18), .E(E_18), .F(F_18), .G(G_18));
	DFSM # (.MAX_nPERIOD(MAX_nPERIOD), .MAX_nLMAC(MAX_nLMAC), .MAX_nSHFT(MAX_nSHFT)) fsm_19(.clk(clk), .rst(rst), .config_en(dfsm_config_en), .iconfig(dfsm_config), .in_en(dfsm_data_en_18), .start(start_bypass_18), .in_en_bypass(dfsm_data_en_19), .out_en(dout_en_19), .start_out(start_bypass_19), .A(A_19), .B(B_19), .C(C_19), .D(D_19), .E(E_19), .F(F_19), .G(G_19));
	DFSM # (.MAX_nPERIOD(MAX_nPERIOD), .MAX_nLMAC(MAX_nLMAC), .MAX_nSHFT(MAX_nSHFT)) fsm_20(.clk(clk), .rst(rst), .config_en(dfsm_config_en), .iconfig(dfsm_config), .in_en(dfsm_data_en_19), .start(start_bypass_19), .in_en_bypass(dfsm_data_en_20), .out_en(dout_en_20), .start_out(start_bypass_20), .A(A_20), .B(B_20), .C(C_20), .D(D_20), .E(E_20), .F(F_20), .G(G_20));
	DFSM # (.MAX_nPERIOD(MAX_nPERIOD), .MAX_nLMAC(MAX_nLMAC), .MAX_nSHFT(MAX_nSHFT)) fsm_21(.clk(clk), .rst(rst), .config_en(dfsm_config_en), .iconfig(dfsm_config), .in_en(dfsm_data_en_20), .start(start_bypass_20), .in_en_bypass(dfsm_data_en_21), .out_en(dout_en_21), .start_out(start_bypass_21), .A(A_21), .B(B_21), .C(C_21), .D(D_21), .E(E_21), .F(F_21), .G(G_21));
	DFSM # (.MAX_nPERIOD(MAX_nPERIOD), .MAX_nLMAC(MAX_nLMAC), .MAX_nSHFT(MAX_nSHFT)) fsm_22(.clk(clk), .rst(rst), .config_en(dfsm_config_en), .iconfig(dfsm_config), .in_en(dfsm_data_en_21), .start(start_bypass_21), .in_en_bypass(dfsm_data_en_22), .out_en(dout_en_22), .start_out(start_bypass_22), .A(A_22), .B(B_22), .C(C_22), .D(D_22), .E(E_22), .F(F_22), .G(G_22));
	DFSM # (.MAX_nPERIOD(MAX_nPERIOD), .MAX_nLMAC(MAX_nLMAC), .MAX_nSHFT(MAX_nSHFT)) fsm_23(.clk(clk), .rst(rst), .config_en(dfsm_config_en), .iconfig(dfsm_config), .in_en(dfsm_data_en_22), .start(start_bypass_22), .in_en_bypass(dfsm_data_en_23), .out_en(dout_en_23), .start_out(start_bypass_23), .A(A_23), .B(B_23), .C(C_23), .D(D_23), .E(E_23), .F(F_23), .G(G_23));
	DFSM # (.MAX_nPERIOD(MAX_nPERIOD), .MAX_nLMAC(MAX_nLMAC), .MAX_nSHFT(MAX_nSHFT)) fsm_24(.clk(clk), .rst(rst), .config_en(dfsm_config_en), .iconfig(dfsm_config), .in_en(dfsm_data_en_23), .start(start_bypass_23), .in_en_bypass(dfsm_data_en_24), .out_en(dout_en_24), .start_out(start_bypass_24), .A(A_24), .B(B_24), .C(C_24), .D(D_24), .E(E_24), .F(F_24), .G(G_24));
	DFSM # (.MAX_nPERIOD(MAX_nPERIOD), .MAX_nLMAC(MAX_nLMAC), .MAX_nSHFT(MAX_nSHFT)) fsm_25(.clk(clk), .rst(rst), .config_en(dfsm_config_en), .iconfig(dfsm_config), .in_en(dfsm_data_en_24), .start(start_bypass_24), .in_en_bypass(dfsm_data_en_25), .out_en(dout_en_25), .start_out(start_bypass_25), .A(A_25), .B(B_25), .C(C_25), .D(D_25), .E(E_25), .F(F_25), .G(G_25));
	DFSM # (.MAX_nPERIOD(MAX_nPERIOD), .MAX_nLMAC(MAX_nLMAC), .MAX_nSHFT(MAX_nSHFT)) fsm_26(.clk(clk), .rst(rst), .config_en(dfsm_config_en), .iconfig(dfsm_config), .in_en(dfsm_data_en_25), .start(start_bypass_25), .in_en_bypass(dfsm_data_en_26), .out_en(dout_en_26), .start_out(start_bypass_26), .A(A_26), .B(B_26), .C(C_26), .D(D_26), .E(E_26), .F(F_26), .G(G_26));
	DFSM # (.MAX_nPERIOD(MAX_nPERIOD), .MAX_nLMAC(MAX_nLMAC), .MAX_nSHFT(MAX_nSHFT)) fsm_27(.clk(clk), .rst(rst), .config_en(dfsm_config_en), .iconfig(dfsm_config), .in_en(dfsm_data_en_26), .start(start_bypass_26), .in_en_bypass(dfsm_data_en_27), .out_en(dout_en_27), .start_out(start_bypass_27), .A(A_27), .B(B_27), .C(C_27), .D(D_27), .E(E_27), .F(F_27), .G(G_27));
	DFSM # (.MAX_nPERIOD(MAX_nPERIOD), .MAX_nLMAC(MAX_nLMAC), .MAX_nSHFT(MAX_nSHFT)) fsm_28(.clk(clk), .rst(rst), .config_en(dfsm_config_en), .iconfig(dfsm_config), .in_en(dfsm_data_en_27), .start(start_bypass_27), .in_en_bypass(dfsm_data_en_28), .out_en(dout_en_28), .start_out(start_bypass_28), .A(A_28), .B(B_28), .C(C_28), .D(D_28), .E(E_28), .F(F_28), .G(G_28));
	DFSM # (.MAX_nPERIOD(MAX_nPERIOD), .MAX_nLMAC(MAX_nLMAC), .MAX_nSHFT(MAX_nSHFT)) fsm_29(.clk(clk), .rst(rst), .config_en(dfsm_config_en), .iconfig(dfsm_config), .in_en(dfsm_data_en_28), .start(start_bypass_28), .in_en_bypass(dfsm_data_en_29), .out_en(dout_en_29), .start_out(start_bypass_29), .A(A_29), .B(B_29), .C(C_29), .D(D_29), .E(E_29), .F(F_29), .G(G_29));
	DFSM # (.MAX_nPERIOD(MAX_nPERIOD), .MAX_nLMAC(MAX_nLMAC), .MAX_nSHFT(MAX_nSHFT)) fsm_30(.clk(clk), .rst(rst), .config_en(dfsm_config_en), .iconfig(dfsm_config), .in_en(dfsm_data_en_29), .start(start_bypass_29), .in_en_bypass(dfsm_data_en_30), .out_en(dout_en_30), .start_out(start_bypass_30), .A(A_30), .B(B_30), .C(C_30), .D(D_30), .E(E_30), .F(F_30), .G(G_30));
	DFSM # (.MAX_nPERIOD(MAX_nPERIOD), .MAX_nLMAC(MAX_nLMAC), .MAX_nSHFT(MAX_nSHFT)) fsm_31(.clk(clk), .rst(rst), .config_en(dfsm_config_en), .iconfig(dfsm_config), .in_en(dfsm_data_en_30), .start(start_bypass_30), .in_en_bypass(dfsm_data_en_31), .out_en(dout_en_31), .start_out(start_bypass_31), .A(A_31), .B(B_31), .C(C_31), .D(D_31), .E(E_31), .F(F_31), .G(G_31));
	DFSM # (.MAX_nPERIOD(MAX_nPERIOD), .MAX_nLMAC(MAX_nLMAC), .MAX_nSHFT(MAX_nSHFT)) fsm_32(.clk(clk), .rst(rst), .config_en(dfsm_config_en), .iconfig(dfsm_config), .in_en(dfsm_data_en_31), .start(start_bypass_31), .in_en_bypass(dfsm_data_en_32), .out_en(dout_en_32), .start_out(start_bypass_32), .A(A_32), .B(B_32), .C(C_32), .D(D_32), .E(E_32), .F(F_32), .G(G_32));

endmodule
