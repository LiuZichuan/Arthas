`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: Liu Zichuan
// 
// Create Date: 09/01/2017 09:40:47 PM
// Design Name: Arthas
// Module Name: SystolicBank
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies:
// 
// Revision: 0.1
// Revision 0.01 - File Created
// Additional Comments:
//
//////////////////////////////////////////////////////////////////////////////////

module SystolicBank(
	// inputs
	clk,
	rst,
	in_en,
	iconfig_1,
	iconfig_2,
	iconfig_3,
	config_load,
	weight_1,
	weight_2,
	weight_3,
	feature_1,
	feature_2,
	feature_3,
	feature_4,
	feature_5,
	feature_6,
	feature_7,
	feature_8,
	feature_9,
	feature_10,
	feature_11,
	feature_12,
	feature_13,
	feature_14,
	feature_15,
	feature_16,
	feature_17,
	feature_18,
	feature_19,
	feature_20,
	feature_21,
	feature_22,
	feature_23,
	feature_24,
	feature_25,
	feature_26,
	feature_27,
	feature_28,
	feature_29,
	feature_30,
	feature_31,
	feature_32,
	feature_33,
	feature_34,
	A_1,
	A_2,
	A_3,
	A_4,
	A_5,
	A_6,
	A_7,
	A_8,
	A_9,
	A_10,
	A_11,
	A_12,
	A_13,
	A_14,
	A_15,
	A_16,
	A_17,
	A_18,
	A_19,
	A_20,
	A_21,
	A_22,
	A_23,
	A_24,
	A_25,
	A_26,
	A_27,
	A_28,
	A_29,
	A_30,
	A_31,
	A_32,
	B_1,
	B_2,
	B_3,
	B_4,
	B_5,
	B_6,
	B_7,
	B_8,
	B_9,
	B_10,
	B_11,
	B_12,
	B_13,
	B_14,
	B_15,
	B_16,
	B_17,
	B_18,
	B_19,
	B_20,
	B_21,
	B_22,
	B_23,
	B_24,
	B_25,
	B_26,
	B_27,
	B_28,
	B_29,
	B_30,
	B_31,
	B_32,
	C_1,
	C_2,
	C_3,
	C_4,
	C_5,
	C_6,
	C_7,
	C_8,
	C_9,
	C_10,
	C_11,
	C_12,
	C_13,
	C_14,
	C_15,
	C_16,
	C_17,
	C_18,
	C_19,
	C_20,
	C_21,
	C_22,
	C_23,
	C_24,
	C_25,
	C_26,
	C_27,
	C_28,
	C_29,
	C_30,
	C_31,
	C_32,
	D_1,
	D_2,
	D_3,
	D_4,
	D_5,
	D_6,
	D_7,
	D_8,
	D_9,
	D_10,
	D_11,
	D_12,
	D_13,
	D_14,
	D_15,
	D_16,
	D_17,
	D_18,
	D_19,
	D_20,
	D_21,
	D_22,
	D_23,
	D_24,
	D_25,
	D_26,
	D_27,
	D_28,
	D_29,
	D_30,
	D_31,
	D_32,
	E_1,
	E_2,
	E_3,
	E_4,
	E_5,
	E_6,
	E_7,
	E_8,
	E_9,
	E_10,
	E_11,
	E_12,
	E_13,
	E_14,
	E_15,
	E_16,
	E_17,
	E_18,
	E_19,
	E_20,
	E_21,
	E_22,
	E_23,
	E_24,
	E_25,
	E_26,
	E_27,
	E_28,
	E_29,
	E_30,
	E_31,
	E_32,
	F_1,
	F_2,
	F_3,
	F_4,
	F_5,
	F_6,
	F_7,
	F_8,
	F_9,
	F_10,
	F_11,
	F_12,
	F_13,
	F_14,
	F_15,
	F_16,
	F_17,
	F_18,
	F_19,
	F_20,
	F_21,
	F_22,
	F_23,
	F_24,
	F_25,
	F_26,
	F_27,
	F_28,
	F_29,
	F_30,
	F_31,
	F_32,
	G_1,
	G_2,
	G_3,
	G_4,
	G_5,
	G_6,
	G_7,
	G_8,
	G_9,
	G_10,
	G_11,
	G_12,
	G_13,
	G_14,
	G_15,
	G_16,
	G_17,
	G_18,
	G_19,
	G_20,
	G_21,
	G_22,
	G_23,
	G_24,
	G_25,
	G_26,
	G_27,
	G_28,
	G_29,
	G_30,
	G_31,
	G_32,
	// outputs
	dout_1,
	dout_2,
	dout_3,
	dout_4,
	dout_5,
	dout_6,
	dout_7,
	dout_8,
	dout_9,
	dout_10,
	dout_11,
	dout_12,
	dout_13,
	dout_14,
	dout_15,
	dout_16,
	dout_17,
	dout_18,
	dout_19,
	dout_20,
	dout_21,
	dout_22,
	dout_23,
	dout_24,
	dout_25,
	dout_26,
	dout_27,
	dout_28,
	dout_29,
	dout_30,
	dout_31,
	dout_32
);
	parameter nCols = 32;
	parameter nRows = 3;
	parameter iWidth = 16;
	parameter oWidth = 33;

	// inputs
	input clk, rst, in_en, config_load;
	input iconfig_1;
	input iconfig_2;
	input iconfig_3;
	input [15:0] weight_1;
	input [15:0] weight_2;
	input [15:0] weight_3;
	input [15:0] feature_1;
	input [15:0] feature_2;
	input [15:0] feature_3;
	input [15:0] feature_4;
	input [15:0] feature_5;
	input [15:0] feature_6;
	input [15:0] feature_7;
	input [15:0] feature_8;
	input [15:0] feature_9;
	input [15:0] feature_10;
	input [15:0] feature_11;
	input [15:0] feature_12;
	input [15:0] feature_13;
	input [15:0] feature_14;
	input [15:0] feature_15;
	input [15:0] feature_16;
	input [15:0] feature_17;
	input [15:0] feature_18;
	input [15:0] feature_19;
	input [15:0] feature_20;
	input [15:0] feature_21;
	input [15:0] feature_22;
	input [15:0] feature_23;
	input [15:0] feature_24;
	input [15:0] feature_25;
	input [15:0] feature_26;
	input [15:0] feature_27;
	input [15:0] feature_28;
	input [15:0] feature_29;
	input [15:0] feature_30;
	input [15:0] feature_31;
	input [15:0] feature_32;
	input [15:0] feature_33;
	input [15:0] feature_34;
	input A_1;
	input A_2;
	input A_3;
	input A_4;
	input A_5;
	input A_6;
	input A_7;
	input A_8;
	input A_9;
	input A_10;
	input A_11;
	input A_12;
	input A_13;
	input A_14;
	input A_15;
	input A_16;
	input A_17;
	input A_18;
	input A_19;
	input A_20;
	input A_21;
	input A_22;
	input A_23;
	input A_24;
	input A_25;
	input A_26;
	input A_27;
	input A_28;
	input A_29;
	input A_30;
	input A_31;
	input A_32;
	input B_1;
	input B_2;
	input B_3;
	input B_4;
	input B_5;
	input B_6;
	input B_7;
	input B_8;
	input B_9;
	input B_10;
	input B_11;
	input B_12;
	input B_13;
	input B_14;
	input B_15;
	input B_16;
	input B_17;
	input B_18;
	input B_19;
	input B_20;
	input B_21;
	input B_22;
	input B_23;
	input B_24;
	input B_25;
	input B_26;
	input B_27;
	input B_28;
	input B_29;
	input B_30;
	input B_31;
	input B_32;
	input C_1;
	input C_2;
	input C_3;
	input C_4;
	input C_5;
	input C_6;
	input C_7;
	input C_8;
	input C_9;
	input C_10;
	input C_11;
	input C_12;
	input C_13;
	input C_14;
	input C_15;
	input C_16;
	input C_17;
	input C_18;
	input C_19;
	input C_20;
	input C_21;
	input C_22;
	input C_23;
	input C_24;
	input C_25;
	input C_26;
	input C_27;
	input C_28;
	input C_29;
	input C_30;
	input C_31;
	input C_32;
	input D_1;
	input D_2;
	input D_3;
	input D_4;
	input D_5;
	input D_6;
	input D_7;
	input D_8;
	input D_9;
	input D_10;
	input D_11;
	input D_12;
	input D_13;
	input D_14;
	input D_15;
	input D_16;
	input D_17;
	input D_18;
	input D_19;
	input D_20;
	input D_21;
	input D_22;
	input D_23;
	input D_24;
	input D_25;
	input D_26;
	input D_27;
	input D_28;
	input D_29;
	input D_30;
	input D_31;
	input D_32;
	input E_1;
	input E_2;
	input E_3;
	input E_4;
	input E_5;
	input E_6;
	input E_7;
	input E_8;
	input E_9;
	input E_10;
	input E_11;
	input E_12;
	input E_13;
	input E_14;
	input E_15;
	input E_16;
	input E_17;
	input E_18;
	input E_19;
	input E_20;
	input E_21;
	input E_22;
	input E_23;
	input E_24;
	input E_25;
	input E_26;
	input E_27;
	input E_28;
	input E_29;
	input E_30;
	input E_31;
	input E_32;
	input F_1;
	input F_2;
	input F_3;
	input F_4;
	input F_5;
	input F_6;
	input F_7;
	input F_8;
	input F_9;
	input F_10;
	input F_11;
	input F_12;
	input F_13;
	input F_14;
	input F_15;
	input F_16;
	input F_17;
	input F_18;
	input F_19;
	input F_20;
	input F_21;
	input F_22;
	input F_23;
	input F_24;
	input F_25;
	input F_26;
	input F_27;
	input F_28;
	input F_29;
	input F_30;
	input F_31;
	input F_32;
	input G_1;
	input G_2;
	input G_3;
	input G_4;
	input G_5;
	input G_6;
	input G_7;
	input G_8;
	input G_9;
	input G_10;
	input G_11;
	input G_12;
	input G_13;
	input G_14;
	input G_15;
	input G_16;
	input G_17;
	input G_18;
	input G_19;
	input G_20;
	input G_21;
	input G_22;
	input G_23;
	input G_24;
	input G_25;
	input G_26;
	input G_27;
	input G_28;
	input G_29;
	input G_30;
	input G_31;
	input G_32;

	// outputs
	output [32:0] dout_1;
	output [32:0] dout_2;
	output [32:0] dout_3;
	output [32:0] dout_4;
	output [32:0] dout_5;
	output [32:0] dout_6;
	output [32:0] dout_7;
	output [32:0] dout_8;
	output [32:0] dout_9;
	output [32:0] dout_10;
	output [32:0] dout_11;
	output [32:0] dout_12;
	output [32:0] dout_13;
	output [32:0] dout_14;
	output [32:0] dout_15;
	output [32:0] dout_16;
	output [32:0] dout_17;
	output [32:0] dout_18;
	output [32:0] dout_19;
	output [32:0] dout_20;
	output [32:0] dout_21;
	output [32:0] dout_22;
	output [32:0] dout_23;
	output [32:0] dout_24;
	output [32:0] dout_25;
	output [32:0] dout_26;
	output [32:0] dout_27;
	output [32:0] dout_28;
	output [32:0] dout_29;
	output [32:0] dout_30;
	output [32:0] dout_31;
	output [32:0] dout_32;

	logic wf_en_1_0;
	logic wf_en_1_1;
	logic wf_en_1_2;
	logic wf_en_1_3;
	logic wf_en_1_4;
	logic wf_en_1_5;
	logic wf_en_1_6;
	logic wf_en_1_7;
	logic wf_en_1_8;
	logic wf_en_1_9;
	logic wf_en_1_10;
	logic wf_en_1_11;
	logic wf_en_1_12;
	logic wf_en_1_13;
	logic wf_en_1_14;
	logic wf_en_1_15;
	logic wf_en_1_16;
	logic wf_en_1_17;
	logic wf_en_1_18;
	logic wf_en_1_19;
	logic wf_en_1_20;
	logic wf_en_1_21;
	logic wf_en_1_22;
	logic wf_en_1_23;
	logic wf_en_1_24;
	logic wf_en_1_25;
	logic wf_en_1_26;
	logic wf_en_1_27;
	logic wf_en_1_28;
	logic wf_en_1_29;
	logic wf_en_1_30;
	logic wf_en_1_31;
	logic wf_en_1_32;
	logic wf_en_2_0;
	logic wf_en_2_1;
	logic wf_en_2_2;
	logic wf_en_2_3;
	logic wf_en_2_4;
	logic wf_en_2_5;
	logic wf_en_2_6;
	logic wf_en_2_7;
	logic wf_en_2_8;
	logic wf_en_2_9;
	logic wf_en_2_10;
	logic wf_en_2_11;
	logic wf_en_2_12;
	logic wf_en_2_13;
	logic wf_en_2_14;
	logic wf_en_2_15;
	logic wf_en_2_16;
	logic wf_en_2_17;
	logic wf_en_2_18;
	logic wf_en_2_19;
	logic wf_en_2_20;
	logic wf_en_2_21;
	logic wf_en_2_22;
	logic wf_en_2_23;
	logic wf_en_2_24;
	logic wf_en_2_25;
	logic wf_en_2_26;
	logic wf_en_2_27;
	logic wf_en_2_28;
	logic wf_en_2_29;
	logic wf_en_2_30;
	logic wf_en_2_31;
	logic wf_en_2_32;
	logic wf_en_3_0;
	logic wf_en_3_1;
	logic wf_en_3_2;
	logic wf_en_3_3;
	logic wf_en_3_4;
	logic wf_en_3_5;
	logic wf_en_3_6;
	logic wf_en_3_7;
	logic wf_en_3_8;
	logic wf_en_3_9;
	logic wf_en_3_10;
	logic wf_en_3_11;
	logic wf_en_3_12;
	logic wf_en_3_13;
	logic wf_en_3_14;
	logic wf_en_3_15;
	logic wf_en_3_16;
	logic wf_en_3_17;
	logic wf_en_3_18;
	logic wf_en_3_19;
	logic wf_en_3_20;
	logic wf_en_3_21;
	logic wf_en_3_22;
	logic wf_en_3_23;
	logic wf_en_3_24;
	logic wf_en_3_25;
	logic wf_en_3_26;
	logic wf_en_3_27;
	logic wf_en_3_28;
	logic wf_en_3_29;
	logic wf_en_3_30;
	logic wf_en_3_31;
	logic wf_en_3_32;

	logic [32:0] psum_1_1;
	logic [32:0] psum_1_2;
	logic [32:0] psum_1_3;
	logic [32:0] psum_1_4;
	logic [32:0] psum_1_5;
	logic [32:0] psum_1_6;
	logic [32:0] psum_1_7;
	logic [32:0] psum_1_8;
	logic [32:0] psum_1_9;
	logic [32:0] psum_1_10;
	logic [32:0] psum_1_11;
	logic [32:0] psum_1_12;
	logic [32:0] psum_1_13;
	logic [32:0] psum_1_14;
	logic [32:0] psum_1_15;
	logic [32:0] psum_1_16;
	logic [32:0] psum_1_17;
	logic [32:0] psum_1_18;
	logic [32:0] psum_1_19;
	logic [32:0] psum_1_20;
	logic [32:0] psum_1_21;
	logic [32:0] psum_1_22;
	logic [32:0] psum_1_23;
	logic [32:0] psum_1_24;
	logic [32:0] psum_1_25;
	logic [32:0] psum_1_26;
	logic [32:0] psum_1_27;
	logic [32:0] psum_1_28;
	logic [32:0] psum_1_29;
	logic [32:0] psum_1_30;
	logic [32:0] psum_1_31;
	logic [32:0] psum_1_32;
	logic [32:0] psum_2_1;
	logic [32:0] psum_2_2;
	logic [32:0] psum_2_3;
	logic [32:0] psum_2_4;
	logic [32:0] psum_2_5;
	logic [32:0] psum_2_6;
	logic [32:0] psum_2_7;
	logic [32:0] psum_2_8;
	logic [32:0] psum_2_9;
	logic [32:0] psum_2_10;
	logic [32:0] psum_2_11;
	logic [32:0] psum_2_12;
	logic [32:0] psum_2_13;
	logic [32:0] psum_2_14;
	logic [32:0] psum_2_15;
	logic [32:0] psum_2_16;
	logic [32:0] psum_2_17;
	logic [32:0] psum_2_18;
	logic [32:0] psum_2_19;
	logic [32:0] psum_2_20;
	logic [32:0] psum_2_21;
	logic [32:0] psum_2_22;
	logic [32:0] psum_2_23;
	logic [32:0] psum_2_24;
	logic [32:0] psum_2_25;
	logic [32:0] psum_2_26;
	logic [32:0] psum_2_27;
	logic [32:0] psum_2_28;
	logic [32:0] psum_2_29;
	logic [32:0] psum_2_30;
	logic [32:0] psum_2_31;
	logic [32:0] psum_2_32;
	logic [32:0] psum_3_1;
	logic [32:0] psum_3_2;
	logic [32:0] psum_3_3;
	logic [32:0] psum_3_4;
	logic [32:0] psum_3_5;
	logic [32:0] psum_3_6;
	logic [32:0] psum_3_7;
	logic [32:0] psum_3_8;
	logic [32:0] psum_3_9;
	logic [32:0] psum_3_10;
	logic [32:0] psum_3_11;
	logic [32:0] psum_3_12;
	logic [32:0] psum_3_13;
	logic [32:0] psum_3_14;
	logic [32:0] psum_3_15;
	logic [32:0] psum_3_16;
	logic [32:0] psum_3_17;
	logic [32:0] psum_3_18;
	logic [32:0] psum_3_19;
	logic [32:0] psum_3_20;
	logic [32:0] psum_3_21;
	logic [32:0] psum_3_22;
	logic [32:0] psum_3_23;
	logic [32:0] psum_3_24;
	logic [32:0] psum_3_25;
	logic [32:0] psum_3_26;
	logic [32:0] psum_3_27;
	logic [32:0] psum_3_28;
	logic [32:0] psum_3_29;
	logic [32:0] psum_3_30;
	logic [32:0] psum_3_31;
	logic [32:0] psum_3_32;
	logic [32:0] psum_4_1;
	logic [32:0] psum_4_2;
	logic [32:0] psum_4_3;
	logic [32:0] psum_4_4;
	logic [32:0] psum_4_5;
	logic [32:0] psum_4_6;
	logic [32:0] psum_4_7;
	logic [32:0] psum_4_8;
	logic [32:0] psum_4_9;
	logic [32:0] psum_4_10;
	logic [32:0] psum_4_11;
	logic [32:0] psum_4_12;
	logic [32:0] psum_4_13;
	logic [32:0] psum_4_14;
	logic [32:0] psum_4_15;
	logic [32:0] psum_4_16;
	logic [32:0] psum_4_17;
	logic [32:0] psum_4_18;
	logic [32:0] psum_4_19;
	logic [32:0] psum_4_20;
	logic [32:0] psum_4_21;
	logic [32:0] psum_4_22;
	logic [32:0] psum_4_23;
	logic [32:0] psum_4_24;
	logic [32:0] psum_4_25;
	logic [32:0] psum_4_26;
	logic [32:0] psum_4_27;
	logic [32:0] psum_4_28;
	logic [32:0] psum_4_29;
	logic [32:0] psum_4_30;
	logic [32:0] psum_4_31;
	logic [32:0] psum_4_32;

	logic [15:0] weight_1_0;
	logic [15:0] weight_1_1;
	logic [15:0] weight_1_2;
	logic [15:0] weight_1_3;
	logic [15:0] weight_1_4;
	logic [15:0] weight_1_5;
	logic [15:0] weight_1_6;
	logic [15:0] weight_1_7;
	logic [15:0] weight_1_8;
	logic [15:0] weight_1_9;
	logic [15:0] weight_1_10;
	logic [15:0] weight_1_11;
	logic [15:0] weight_1_12;
	logic [15:0] weight_1_13;
	logic [15:0] weight_1_14;
	logic [15:0] weight_1_15;
	logic [15:0] weight_1_16;
	logic [15:0] weight_1_17;
	logic [15:0] weight_1_18;
	logic [15:0] weight_1_19;
	logic [15:0] weight_1_20;
	logic [15:0] weight_1_21;
	logic [15:0] weight_1_22;
	logic [15:0] weight_1_23;
	logic [15:0] weight_1_24;
	logic [15:0] weight_1_25;
	logic [15:0] weight_1_26;
	logic [15:0] weight_1_27;
	logic [15:0] weight_1_28;
	logic [15:0] weight_1_29;
	logic [15:0] weight_1_30;
	logic [15:0] weight_1_31;
	logic [15:0] weight_1_32;
	logic [15:0] weight_2_0;
	logic [15:0] weight_2_1;
	logic [15:0] weight_2_2;
	logic [15:0] weight_2_3;
	logic [15:0] weight_2_4;
	logic [15:0] weight_2_5;
	logic [15:0] weight_2_6;
	logic [15:0] weight_2_7;
	logic [15:0] weight_2_8;
	logic [15:0] weight_2_9;
	logic [15:0] weight_2_10;
	logic [15:0] weight_2_11;
	logic [15:0] weight_2_12;
	logic [15:0] weight_2_13;
	logic [15:0] weight_2_14;
	logic [15:0] weight_2_15;
	logic [15:0] weight_2_16;
	logic [15:0] weight_2_17;
	logic [15:0] weight_2_18;
	logic [15:0] weight_2_19;
	logic [15:0] weight_2_20;
	logic [15:0] weight_2_21;
	logic [15:0] weight_2_22;
	logic [15:0] weight_2_23;
	logic [15:0] weight_2_24;
	logic [15:0] weight_2_25;
	logic [15:0] weight_2_26;
	logic [15:0] weight_2_27;
	logic [15:0] weight_2_28;
	logic [15:0] weight_2_29;
	logic [15:0] weight_2_30;
	logic [15:0] weight_2_31;
	logic [15:0] weight_2_32;
	logic [15:0] weight_3_0;
	logic [15:0] weight_3_1;
	logic [15:0] weight_3_2;
	logic [15:0] weight_3_3;
	logic [15:0] weight_3_4;
	logic [15:0] weight_3_5;
	logic [15:0] weight_3_6;
	logic [15:0] weight_3_7;
	logic [15:0] weight_3_8;
	logic [15:0] weight_3_9;
	logic [15:0] weight_3_10;
	logic [15:0] weight_3_11;
	logic [15:0] weight_3_12;
	logic [15:0] weight_3_13;
	logic [15:0] weight_3_14;
	logic [15:0] weight_3_15;
	logic [15:0] weight_3_16;
	logic [15:0] weight_3_17;
	logic [15:0] weight_3_18;
	logic [15:0] weight_3_19;
	logic [15:0] weight_3_20;
	logic [15:0] weight_3_21;
	logic [15:0] weight_3_22;
	logic [15:0] weight_3_23;
	logic [15:0] weight_3_24;
	logic [15:0] weight_3_25;
	logic [15:0] weight_3_26;
	logic [15:0] weight_3_27;
	logic [15:0] weight_3_28;
	logic [15:0] weight_3_29;
	logic [15:0] weight_3_30;
	logic [15:0] weight_3_31;
	logic [15:0] weight_3_32;
	logic [15:0] weight_4_0;
	logic [15:0] weight_4_1;
	logic [15:0] weight_4_2;
	logic [15:0] weight_4_3;
	logic [15:0] weight_4_4;
	logic [15:0] weight_4_5;
	logic [15:0] weight_4_6;
	logic [15:0] weight_4_7;
	logic [15:0] weight_4_8;
	logic [15:0] weight_4_9;
	logic [15:0] weight_4_10;
	logic [15:0] weight_4_11;
	logic [15:0] weight_4_12;
	logic [15:0] weight_4_13;
	logic [15:0] weight_4_14;
	logic [15:0] weight_4_15;
	logic [15:0] weight_4_16;
	logic [15:0] weight_4_17;
	logic [15:0] weight_4_18;
	logic [15:0] weight_4_19;
	logic [15:0] weight_4_20;
	logic [15:0] weight_4_21;
	logic [15:0] weight_4_22;
	logic [15:0] weight_4_23;
	logic [15:0] weight_4_24;
	logic [15:0] weight_4_25;
	logic [15:0] weight_4_26;
	logic [15:0] weight_4_27;
	logic [15:0] weight_4_28;
	logic [15:0] weight_4_29;
	logic [15:0] weight_4_30;
	logic [15:0] weight_4_31;
	logic [15:0] weight_4_32;

	logic [15:0] feature_1_0;
	logic [15:0] feature_1_1;
	logic [15:0] feature_1_2;
	logic [15:0] feature_1_3;
	logic [15:0] feature_1_4;
	logic [15:0] feature_1_5;
	logic [15:0] feature_1_6;
	logic [15:0] feature_1_7;
	logic [15:0] feature_1_8;
	logic [15:0] feature_1_9;
	logic [15:0] feature_1_10;
	logic [15:0] feature_1_11;
	logic [15:0] feature_1_12;
	logic [15:0] feature_1_13;
	logic [15:0] feature_1_14;
	logic [15:0] feature_1_15;
	logic [15:0] feature_1_16;
	logic [15:0] feature_1_17;
	logic [15:0] feature_1_18;
	logic [15:0] feature_1_19;
	logic [15:0] feature_1_20;
	logic [15:0] feature_1_21;
	logic [15:0] feature_1_22;
	logic [15:0] feature_1_23;
	logic [15:0] feature_1_24;
	logic [15:0] feature_1_25;
	logic [15:0] feature_1_26;
	logic [15:0] feature_1_27;
	logic [15:0] feature_1_28;
	logic [15:0] feature_1_29;
	logic [15:0] feature_1_30;
	logic [15:0] feature_1_31;
	logic [15:0] feature_1_32;
	logic [15:0] feature_2_0;
	logic [15:0] feature_2_1;
	logic [15:0] feature_2_2;
	logic [15:0] feature_2_3;
	logic [15:0] feature_2_4;
	logic [15:0] feature_2_5;
	logic [15:0] feature_2_6;
	logic [15:0] feature_2_7;
	logic [15:0] feature_2_8;
	logic [15:0] feature_2_9;
	logic [15:0] feature_2_10;
	logic [15:0] feature_2_11;
	logic [15:0] feature_2_12;
	logic [15:0] feature_2_13;
	logic [15:0] feature_2_14;
	logic [15:0] feature_2_15;
	logic [15:0] feature_2_16;
	logic [15:0] feature_2_17;
	logic [15:0] feature_2_18;
	logic [15:0] feature_2_19;
	logic [15:0] feature_2_20;
	logic [15:0] feature_2_21;
	logic [15:0] feature_2_22;
	logic [15:0] feature_2_23;
	logic [15:0] feature_2_24;
	logic [15:0] feature_2_25;
	logic [15:0] feature_2_26;
	logic [15:0] feature_2_27;
	logic [15:0] feature_2_28;
	logic [15:0] feature_2_29;
	logic [15:0] feature_2_30;
	logic [15:0] feature_2_31;
	logic [15:0] feature_2_32;
	logic [15:0] feature_3_0;
	logic [15:0] feature_3_1;
	logic [15:0] feature_3_2;
	logic [15:0] feature_3_3;
	logic [15:0] feature_3_4;
	logic [15:0] feature_3_5;
	logic [15:0] feature_3_6;
	logic [15:0] feature_3_7;
	logic [15:0] feature_3_8;
	logic [15:0] feature_3_9;
	logic [15:0] feature_3_10;
	logic [15:0] feature_3_11;
	logic [15:0] feature_3_12;
	logic [15:0] feature_3_13;
	logic [15:0] feature_3_14;
	logic [15:0] feature_3_15;
	logic [15:0] feature_3_16;
	logic [15:0] feature_3_17;
	logic [15:0] feature_3_18;
	logic [15:0] feature_3_19;
	logic [15:0] feature_3_20;
	logic [15:0] feature_3_21;
	logic [15:0] feature_3_22;
	logic [15:0] feature_3_23;
	logic [15:0] feature_3_24;
	logic [15:0] feature_3_25;
	logic [15:0] feature_3_26;
	logic [15:0] feature_3_27;
	logic [15:0] feature_3_28;
	logic [15:0] feature_3_29;
	logic [15:0] feature_3_30;
	logic [15:0] feature_3_31;
	logic [15:0] feature_3_32;
	logic [15:0] feature_4_0;
	logic [15:0] feature_4_1;
	logic [15:0] feature_4_2;
	logic [15:0] feature_4_3;
	logic [15:0] feature_4_4;
	logic [15:0] feature_4_5;
	logic [15:0] feature_4_6;
	logic [15:0] feature_4_7;
	logic [15:0] feature_4_8;
	logic [15:0] feature_4_9;
	logic [15:0] feature_4_10;
	logic [15:0] feature_4_11;
	logic [15:0] feature_4_12;
	logic [15:0] feature_4_13;
	logic [15:0] feature_4_14;
	logic [15:0] feature_4_15;
	logic [15:0] feature_4_16;
	logic [15:0] feature_4_17;
	logic [15:0] feature_4_18;
	logic [15:0] feature_4_19;
	logic [15:0] feature_4_20;
	logic [15:0] feature_4_21;
	logic [15:0] feature_4_22;
	logic [15:0] feature_4_23;
	logic [15:0] feature_4_24;
	logic [15:0] feature_4_25;
	logic [15:0] feature_4_26;
	logic [15:0] feature_4_27;
	logic [15:0] feature_4_28;
	logic [15:0] feature_4_29;
	logic [15:0] feature_4_30;
	logic [15:0] feature_4_31;
	logic [15:0] feature_4_32;

	assign psum_4_1 = 0;
	assign psum_4_2 = 0;
	assign psum_4_3 = 0;
	assign psum_4_4 = 0;
	assign psum_4_5 = 0;
	assign psum_4_6 = 0;
	assign psum_4_7 = 0;
	assign psum_4_8 = 0;
	assign psum_4_9 = 0;
	assign psum_4_10 = 0;
	assign psum_4_11 = 0;
	assign psum_4_12 = 0;
	assign psum_4_13 = 0;
	assign psum_4_14 = 0;
	assign psum_4_15 = 0;
	assign psum_4_16 = 0;
	assign psum_4_17 = 0;
	assign psum_4_18 = 0;
	assign psum_4_19 = 0;
	assign psum_4_20 = 0;
	assign psum_4_21 = 0;
	assign psum_4_22 = 0;
	assign psum_4_23 = 0;
	assign psum_4_24 = 0;
	assign psum_4_25 = 0;
	assign psum_4_26 = 0;
	assign psum_4_27 = 0;
	assign psum_4_28 = 0;
	assign psum_4_29 = 0;
	assign psum_4_30 = 0;
	assign psum_4_31 = 0;
	assign psum_4_32 = 0;

	assign wf_en_1_0 = in_en;
	assign wf_en_2_0 = in_en;
	assign wf_en_3_0 = in_en;

	assign weight_1_0 = weight_1;
	assign weight_2_0 = weight_2;
	assign weight_3_0 = weight_3;

	assign feature_2_0 = feature_1;
	assign feature_3_0 = feature_2;
	assign feature_4_0 = feature_3;
	assign feature_4_1 = feature_4;
	assign feature_4_2 = feature_5;
	assign feature_4_3 = feature_6;
	assign feature_4_4 = feature_7;
	assign feature_4_5 = feature_8;
	assign feature_4_6 = feature_9;
	assign feature_4_7 = feature_10;
	assign feature_4_8 = feature_11;
	assign feature_4_9 = feature_12;
	assign feature_4_10 = feature_13;
	assign feature_4_11 = feature_14;
	assign feature_4_12 = feature_15;
	assign feature_4_13 = feature_16;
	assign feature_4_14 = feature_17;
	assign feature_4_15 = feature_18;
	assign feature_4_16 = feature_19;
	assign feature_4_17 = feature_20;
	assign feature_4_18 = feature_21;
	assign feature_4_19 = feature_22;
	assign feature_4_20 = feature_23;
	assign feature_4_21 = feature_24;
	assign feature_4_22 = feature_25;
	assign feature_4_23 = feature_26;
	assign feature_4_24 = feature_27;
	assign feature_4_25 = feature_28;
	assign feature_4_26 = feature_29;
	assign feature_4_27 = feature_30;
	assign feature_4_28 = feature_31;
	assign feature_4_29 = feature_32;
	assign feature_4_30 = feature_33;
	assign feature_4_31 = feature_34;

	PEv2 # (.WIDTH(iWidth)) p_1_1(.clk(clk), .rst(rst), .in_en(wf_en_1_0), .ipsum(psum_2_1), .iconfig(iconfig_1), .weight(weight_1_0), .feature(feature_2_0), .config_load(config_load), .A(A_1), .B(B_1), .C(C_1), .D(D_1), .E(E_1), .w_out(weight_1_1), .f_out(feature_1_1), .wf_en(wf_en_1_1), .opsum(psum_1_1));
	PEv2 # (.WIDTH(iWidth)) p_1_2(.clk(clk), .rst(rst), .in_en(wf_en_1_1), .ipsum(psum_2_2), .iconfig(iconfig_1), .weight(weight_1_1), .feature(feature_2_1), .config_load(config_load), .A(A_2), .B(B_2), .C(C_2), .D(D_2), .E(E_2), .w_out(weight_1_2), .f_out(feature_1_2), .wf_en(wf_en_1_2), .opsum(psum_1_2));
	PEv2 # (.WIDTH(iWidth)) p_1_3(.clk(clk), .rst(rst), .in_en(wf_en_1_2), .ipsum(psum_2_3), .iconfig(iconfig_1), .weight(weight_1_2), .feature(feature_2_2), .config_load(config_load), .A(A_3), .B(B_3), .C(C_3), .D(D_3), .E(E_3), .w_out(weight_1_3), .f_out(feature_1_3), .wf_en(wf_en_1_3), .opsum(psum_1_3));
	PEv2 # (.WIDTH(iWidth)) p_1_4(.clk(clk), .rst(rst), .in_en(wf_en_1_3), .ipsum(psum_2_4), .iconfig(iconfig_1), .weight(weight_1_3), .feature(feature_2_3), .config_load(config_load), .A(A_4), .B(B_4), .C(C_4), .D(D_4), .E(E_4), .w_out(weight_1_4), .f_out(feature_1_4), .wf_en(wf_en_1_4), .opsum(psum_1_4));
	PEv2 # (.WIDTH(iWidth)) p_1_5(.clk(clk), .rst(rst), .in_en(wf_en_1_4), .ipsum(psum_2_5), .iconfig(iconfig_1), .weight(weight_1_4), .feature(feature_2_4), .config_load(config_load), .A(A_5), .B(B_5), .C(C_5), .D(D_5), .E(E_5), .w_out(weight_1_5), .f_out(feature_1_5), .wf_en(wf_en_1_5), .opsum(psum_1_5));
	PEv2 # (.WIDTH(iWidth)) p_1_6(.clk(clk), .rst(rst), .in_en(wf_en_1_5), .ipsum(psum_2_6), .iconfig(iconfig_1), .weight(weight_1_5), .feature(feature_2_5), .config_load(config_load), .A(A_6), .B(B_6), .C(C_6), .D(D_6), .E(E_6), .w_out(weight_1_6), .f_out(feature_1_6), .wf_en(wf_en_1_6), .opsum(psum_1_6));
	PEv2 # (.WIDTH(iWidth)) p_1_7(.clk(clk), .rst(rst), .in_en(wf_en_1_6), .ipsum(psum_2_7), .iconfig(iconfig_1), .weight(weight_1_6), .feature(feature_2_6), .config_load(config_load), .A(A_7), .B(B_7), .C(C_7), .D(D_7), .E(E_7), .w_out(weight_1_7), .f_out(feature_1_7), .wf_en(wf_en_1_7), .opsum(psum_1_7));
	PEv2 # (.WIDTH(iWidth)) p_1_8(.clk(clk), .rst(rst), .in_en(wf_en_1_7), .ipsum(psum_2_8), .iconfig(iconfig_1), .weight(weight_1_7), .feature(feature_2_7), .config_load(config_load), .A(A_8), .B(B_8), .C(C_8), .D(D_8), .E(E_8), .w_out(weight_1_8), .f_out(feature_1_8), .wf_en(wf_en_1_8), .opsum(psum_1_8));
	PEv2 # (.WIDTH(iWidth)) p_1_9(.clk(clk), .rst(rst), .in_en(wf_en_1_8), .ipsum(psum_2_9), .iconfig(iconfig_1), .weight(weight_1_8), .feature(feature_2_8), .config_load(config_load), .A(A_9), .B(B_9), .C(C_9), .D(D_9), .E(E_9), .w_out(weight_1_9), .f_out(feature_1_9), .wf_en(wf_en_1_9), .opsum(psum_1_9));
	PEv2 # (.WIDTH(iWidth)) p_1_10(.clk(clk), .rst(rst), .in_en(wf_en_1_9), .ipsum(psum_2_10), .iconfig(iconfig_1), .weight(weight_1_9), .feature(feature_2_9), .config_load(config_load), .A(A_10), .B(B_10), .C(C_10), .D(D_10), .E(E_10), .w_out(weight_1_10), .f_out(feature_1_10), .wf_en(wf_en_1_10), .opsum(psum_1_10));
	PEv2 # (.WIDTH(iWidth)) p_1_11(.clk(clk), .rst(rst), .in_en(wf_en_1_10), .ipsum(psum_2_11), .iconfig(iconfig_1), .weight(weight_1_10), .feature(feature_2_10), .config_load(config_load), .A(A_11), .B(B_11), .C(C_11), .D(D_11), .E(E_11), .w_out(weight_1_11), .f_out(feature_1_11), .wf_en(wf_en_1_11), .opsum(psum_1_11));
	PEv2 # (.WIDTH(iWidth)) p_1_12(.clk(clk), .rst(rst), .in_en(wf_en_1_11), .ipsum(psum_2_12), .iconfig(iconfig_1), .weight(weight_1_11), .feature(feature_2_11), .config_load(config_load), .A(A_12), .B(B_12), .C(C_12), .D(D_12), .E(E_12), .w_out(weight_1_12), .f_out(feature_1_12), .wf_en(wf_en_1_12), .opsum(psum_1_12));
	PEv2 # (.WIDTH(iWidth)) p_1_13(.clk(clk), .rst(rst), .in_en(wf_en_1_12), .ipsum(psum_2_13), .iconfig(iconfig_1), .weight(weight_1_12), .feature(feature_2_12), .config_load(config_load), .A(A_13), .B(B_13), .C(C_13), .D(D_13), .E(E_13), .w_out(weight_1_13), .f_out(feature_1_13), .wf_en(wf_en_1_13), .opsum(psum_1_13));
	PEv2 # (.WIDTH(iWidth)) p_1_14(.clk(clk), .rst(rst), .in_en(wf_en_1_13), .ipsum(psum_2_14), .iconfig(iconfig_1), .weight(weight_1_13), .feature(feature_2_13), .config_load(config_load), .A(A_14), .B(B_14), .C(C_14), .D(D_14), .E(E_14), .w_out(weight_1_14), .f_out(feature_1_14), .wf_en(wf_en_1_14), .opsum(psum_1_14));
	PEv2 # (.WIDTH(iWidth)) p_1_15(.clk(clk), .rst(rst), .in_en(wf_en_1_14), .ipsum(psum_2_15), .iconfig(iconfig_1), .weight(weight_1_14), .feature(feature_2_14), .config_load(config_load), .A(A_15), .B(B_15), .C(C_15), .D(D_15), .E(E_15), .w_out(weight_1_15), .f_out(feature_1_15), .wf_en(wf_en_1_15), .opsum(psum_1_15));
	PEv2 # (.WIDTH(iWidth)) p_1_16(.clk(clk), .rst(rst), .in_en(wf_en_1_15), .ipsum(psum_2_16), .iconfig(iconfig_1), .weight(weight_1_15), .feature(feature_2_15), .config_load(config_load), .A(A_16), .B(B_16), .C(C_16), .D(D_16), .E(E_16), .w_out(weight_1_16), .f_out(feature_1_16), .wf_en(wf_en_1_16), .opsum(psum_1_16));
	PEv2 # (.WIDTH(iWidth)) p_1_17(.clk(clk), .rst(rst), .in_en(wf_en_1_16), .ipsum(psum_2_17), .iconfig(iconfig_1), .weight(weight_1_16), .feature(feature_2_16), .config_load(config_load), .A(A_17), .B(B_17), .C(C_17), .D(D_17), .E(E_17), .w_out(weight_1_17), .f_out(feature_1_17), .wf_en(wf_en_1_17), .opsum(psum_1_17));
	PEv2 # (.WIDTH(iWidth)) p_1_18(.clk(clk), .rst(rst), .in_en(wf_en_1_17), .ipsum(psum_2_18), .iconfig(iconfig_1), .weight(weight_1_17), .feature(feature_2_17), .config_load(config_load), .A(A_18), .B(B_18), .C(C_18), .D(D_18), .E(E_18), .w_out(weight_1_18), .f_out(feature_1_18), .wf_en(wf_en_1_18), .opsum(psum_1_18));
	PEv2 # (.WIDTH(iWidth)) p_1_19(.clk(clk), .rst(rst), .in_en(wf_en_1_18), .ipsum(psum_2_19), .iconfig(iconfig_1), .weight(weight_1_18), .feature(feature_2_18), .config_load(config_load), .A(A_19), .B(B_19), .C(C_19), .D(D_19), .E(E_19), .w_out(weight_1_19), .f_out(feature_1_19), .wf_en(wf_en_1_19), .opsum(psum_1_19));
	PEv2 # (.WIDTH(iWidth)) p_1_20(.clk(clk), .rst(rst), .in_en(wf_en_1_19), .ipsum(psum_2_20), .iconfig(iconfig_1), .weight(weight_1_19), .feature(feature_2_19), .config_load(config_load), .A(A_20), .B(B_20), .C(C_20), .D(D_20), .E(E_20), .w_out(weight_1_20), .f_out(feature_1_20), .wf_en(wf_en_1_20), .opsum(psum_1_20));
	PEv2 # (.WIDTH(iWidth)) p_1_21(.clk(clk), .rst(rst), .in_en(wf_en_1_20), .ipsum(psum_2_21), .iconfig(iconfig_1), .weight(weight_1_20), .feature(feature_2_20), .config_load(config_load), .A(A_21), .B(B_21), .C(C_21), .D(D_21), .E(E_21), .w_out(weight_1_21), .f_out(feature_1_21), .wf_en(wf_en_1_21), .opsum(psum_1_21));
	PEv2 # (.WIDTH(iWidth)) p_1_22(.clk(clk), .rst(rst), .in_en(wf_en_1_21), .ipsum(psum_2_22), .iconfig(iconfig_1), .weight(weight_1_21), .feature(feature_2_21), .config_load(config_load), .A(A_22), .B(B_22), .C(C_22), .D(D_22), .E(E_22), .w_out(weight_1_22), .f_out(feature_1_22), .wf_en(wf_en_1_22), .opsum(psum_1_22));
	PEv2 # (.WIDTH(iWidth)) p_1_23(.clk(clk), .rst(rst), .in_en(wf_en_1_22), .ipsum(psum_2_23), .iconfig(iconfig_1), .weight(weight_1_22), .feature(feature_2_22), .config_load(config_load), .A(A_23), .B(B_23), .C(C_23), .D(D_23), .E(E_23), .w_out(weight_1_23), .f_out(feature_1_23), .wf_en(wf_en_1_23), .opsum(psum_1_23));
	PEv2 # (.WIDTH(iWidth)) p_1_24(.clk(clk), .rst(rst), .in_en(wf_en_1_23), .ipsum(psum_2_24), .iconfig(iconfig_1), .weight(weight_1_23), .feature(feature_2_23), .config_load(config_load), .A(A_24), .B(B_24), .C(C_24), .D(D_24), .E(E_24), .w_out(weight_1_24), .f_out(feature_1_24), .wf_en(wf_en_1_24), .opsum(psum_1_24));
	PEv2 # (.WIDTH(iWidth)) p_1_25(.clk(clk), .rst(rst), .in_en(wf_en_1_24), .ipsum(psum_2_25), .iconfig(iconfig_1), .weight(weight_1_24), .feature(feature_2_24), .config_load(config_load), .A(A_25), .B(B_25), .C(C_25), .D(D_25), .E(E_25), .w_out(weight_1_25), .f_out(feature_1_25), .wf_en(wf_en_1_25), .opsum(psum_1_25));
	PEv2 # (.WIDTH(iWidth)) p_1_26(.clk(clk), .rst(rst), .in_en(wf_en_1_25), .ipsum(psum_2_26), .iconfig(iconfig_1), .weight(weight_1_25), .feature(feature_2_25), .config_load(config_load), .A(A_26), .B(B_26), .C(C_26), .D(D_26), .E(E_26), .w_out(weight_1_26), .f_out(feature_1_26), .wf_en(wf_en_1_26), .opsum(psum_1_26));
	PEv2 # (.WIDTH(iWidth)) p_1_27(.clk(clk), .rst(rst), .in_en(wf_en_1_26), .ipsum(psum_2_27), .iconfig(iconfig_1), .weight(weight_1_26), .feature(feature_2_26), .config_load(config_load), .A(A_27), .B(B_27), .C(C_27), .D(D_27), .E(E_27), .w_out(weight_1_27), .f_out(feature_1_27), .wf_en(wf_en_1_27), .opsum(psum_1_27));
	PEv2 # (.WIDTH(iWidth)) p_1_28(.clk(clk), .rst(rst), .in_en(wf_en_1_27), .ipsum(psum_2_28), .iconfig(iconfig_1), .weight(weight_1_27), .feature(feature_2_27), .config_load(config_load), .A(A_28), .B(B_28), .C(C_28), .D(D_28), .E(E_28), .w_out(weight_1_28), .f_out(feature_1_28), .wf_en(wf_en_1_28), .opsum(psum_1_28));
	PEv2 # (.WIDTH(iWidth)) p_1_29(.clk(clk), .rst(rst), .in_en(wf_en_1_28), .ipsum(psum_2_29), .iconfig(iconfig_1), .weight(weight_1_28), .feature(feature_2_28), .config_load(config_load), .A(A_29), .B(B_29), .C(C_29), .D(D_29), .E(E_29), .w_out(weight_1_29), .f_out(feature_1_29), .wf_en(wf_en_1_29), .opsum(psum_1_29));
	PEv2 # (.WIDTH(iWidth)) p_1_30(.clk(clk), .rst(rst), .in_en(wf_en_1_29), .ipsum(psum_2_30), .iconfig(iconfig_1), .weight(weight_1_29), .feature(feature_2_29), .config_load(config_load), .A(A_30), .B(B_30), .C(C_30), .D(D_30), .E(E_30), .w_out(weight_1_30), .f_out(feature_1_30), .wf_en(wf_en_1_30), .opsum(psum_1_30));
	PEv2 # (.WIDTH(iWidth)) p_1_31(.clk(clk), .rst(rst), .in_en(wf_en_1_30), .ipsum(psum_2_31), .iconfig(iconfig_1), .weight(weight_1_30), .feature(feature_2_30), .config_load(config_load), .A(A_31), .B(B_31), .C(C_31), .D(D_31), .E(E_31), .w_out(weight_1_31), .f_out(feature_1_31), .wf_en(wf_en_1_31), .opsum(psum_1_31));
	PEv2 # (.WIDTH(iWidth)) p_1_32(.clk(clk), .rst(rst), .in_en(wf_en_1_31), .ipsum(psum_2_32), .iconfig(iconfig_1), .weight(weight_1_31), .feature(feature_2_31), .config_load(config_load), .A(A_32), .B(B_32), .C(C_32), .D(D_32), .E(E_32), .w_out(weight_1_32), .f_out(feature_1_32), .wf_en(wf_en_1_32), .opsum(psum_1_32));
	PEv2 # (.WIDTH(iWidth)) p_2_1(.clk(clk), .rst(rst), .in_en(wf_en_2_0), .ipsum(psum_3_1), .iconfig(iconfig_2), .weight(weight_2_0), .feature(feature_3_0), .config_load(config_load), .A(A_1), .B(B_1), .C(C_1), .D(D_1), .E(E_1), .w_out(weight_2_1), .f_out(feature_2_1), .wf_en(wf_en_2_1), .opsum(psum_2_1));
	PEv2 # (.WIDTH(iWidth)) p_2_2(.clk(clk), .rst(rst), .in_en(wf_en_2_1), .ipsum(psum_3_2), .iconfig(iconfig_2), .weight(weight_2_1), .feature(feature_3_1), .config_load(config_load), .A(A_2), .B(B_2), .C(C_2), .D(D_2), .E(E_2), .w_out(weight_2_2), .f_out(feature_2_2), .wf_en(wf_en_2_2), .opsum(psum_2_2));
	PEv2 # (.WIDTH(iWidth)) p_2_3(.clk(clk), .rst(rst), .in_en(wf_en_2_2), .ipsum(psum_3_3), .iconfig(iconfig_2), .weight(weight_2_2), .feature(feature_3_2), .config_load(config_load), .A(A_3), .B(B_3), .C(C_3), .D(D_3), .E(E_3), .w_out(weight_2_3), .f_out(feature_2_3), .wf_en(wf_en_2_3), .opsum(psum_2_3));
	PEv2 # (.WIDTH(iWidth)) p_2_4(.clk(clk), .rst(rst), .in_en(wf_en_2_3), .ipsum(psum_3_4), .iconfig(iconfig_2), .weight(weight_2_3), .feature(feature_3_3), .config_load(config_load), .A(A_4), .B(B_4), .C(C_4), .D(D_4), .E(E_4), .w_out(weight_2_4), .f_out(feature_2_4), .wf_en(wf_en_2_4), .opsum(psum_2_4));
	PEv2 # (.WIDTH(iWidth)) p_2_5(.clk(clk), .rst(rst), .in_en(wf_en_2_4), .ipsum(psum_3_5), .iconfig(iconfig_2), .weight(weight_2_4), .feature(feature_3_4), .config_load(config_load), .A(A_5), .B(B_5), .C(C_5), .D(D_5), .E(E_5), .w_out(weight_2_5), .f_out(feature_2_5), .wf_en(wf_en_2_5), .opsum(psum_2_5));
	PEv2 # (.WIDTH(iWidth)) p_2_6(.clk(clk), .rst(rst), .in_en(wf_en_2_5), .ipsum(psum_3_6), .iconfig(iconfig_2), .weight(weight_2_5), .feature(feature_3_5), .config_load(config_load), .A(A_6), .B(B_6), .C(C_6), .D(D_6), .E(E_6), .w_out(weight_2_6), .f_out(feature_2_6), .wf_en(wf_en_2_6), .opsum(psum_2_6));
	PEv2 # (.WIDTH(iWidth)) p_2_7(.clk(clk), .rst(rst), .in_en(wf_en_2_6), .ipsum(psum_3_7), .iconfig(iconfig_2), .weight(weight_2_6), .feature(feature_3_6), .config_load(config_load), .A(A_7), .B(B_7), .C(C_7), .D(D_7), .E(E_7), .w_out(weight_2_7), .f_out(feature_2_7), .wf_en(wf_en_2_7), .opsum(psum_2_7));
	PEv2 # (.WIDTH(iWidth)) p_2_8(.clk(clk), .rst(rst), .in_en(wf_en_2_7), .ipsum(psum_3_8), .iconfig(iconfig_2), .weight(weight_2_7), .feature(feature_3_7), .config_load(config_load), .A(A_8), .B(B_8), .C(C_8), .D(D_8), .E(E_8), .w_out(weight_2_8), .f_out(feature_2_8), .wf_en(wf_en_2_8), .opsum(psum_2_8));
	PEv2 # (.WIDTH(iWidth)) p_2_9(.clk(clk), .rst(rst), .in_en(wf_en_2_8), .ipsum(psum_3_9), .iconfig(iconfig_2), .weight(weight_2_8), .feature(feature_3_8), .config_load(config_load), .A(A_9), .B(B_9), .C(C_9), .D(D_9), .E(E_9), .w_out(weight_2_9), .f_out(feature_2_9), .wf_en(wf_en_2_9), .opsum(psum_2_9));
	PEv2 # (.WIDTH(iWidth)) p_2_10(.clk(clk), .rst(rst), .in_en(wf_en_2_9), .ipsum(psum_3_10), .iconfig(iconfig_2), .weight(weight_2_9), .feature(feature_3_9), .config_load(config_load), .A(A_10), .B(B_10), .C(C_10), .D(D_10), .E(E_10), .w_out(weight_2_10), .f_out(feature_2_10), .wf_en(wf_en_2_10), .opsum(psum_2_10));
	PEv2 # (.WIDTH(iWidth)) p_2_11(.clk(clk), .rst(rst), .in_en(wf_en_2_10), .ipsum(psum_3_11), .iconfig(iconfig_2), .weight(weight_2_10), .feature(feature_3_10), .config_load(config_load), .A(A_11), .B(B_11), .C(C_11), .D(D_11), .E(E_11), .w_out(weight_2_11), .f_out(feature_2_11), .wf_en(wf_en_2_11), .opsum(psum_2_11));
	PEv2 # (.WIDTH(iWidth)) p_2_12(.clk(clk), .rst(rst), .in_en(wf_en_2_11), .ipsum(psum_3_12), .iconfig(iconfig_2), .weight(weight_2_11), .feature(feature_3_11), .config_load(config_load), .A(A_12), .B(B_12), .C(C_12), .D(D_12), .E(E_12), .w_out(weight_2_12), .f_out(feature_2_12), .wf_en(wf_en_2_12), .opsum(psum_2_12));
	PEv2 # (.WIDTH(iWidth)) p_2_13(.clk(clk), .rst(rst), .in_en(wf_en_2_12), .ipsum(psum_3_13), .iconfig(iconfig_2), .weight(weight_2_12), .feature(feature_3_12), .config_load(config_load), .A(A_13), .B(B_13), .C(C_13), .D(D_13), .E(E_13), .w_out(weight_2_13), .f_out(feature_2_13), .wf_en(wf_en_2_13), .opsum(psum_2_13));
	PEv2 # (.WIDTH(iWidth)) p_2_14(.clk(clk), .rst(rst), .in_en(wf_en_2_13), .ipsum(psum_3_14), .iconfig(iconfig_2), .weight(weight_2_13), .feature(feature_3_13), .config_load(config_load), .A(A_14), .B(B_14), .C(C_14), .D(D_14), .E(E_14), .w_out(weight_2_14), .f_out(feature_2_14), .wf_en(wf_en_2_14), .opsum(psum_2_14));
	PEv2 # (.WIDTH(iWidth)) p_2_15(.clk(clk), .rst(rst), .in_en(wf_en_2_14), .ipsum(psum_3_15), .iconfig(iconfig_2), .weight(weight_2_14), .feature(feature_3_14), .config_load(config_load), .A(A_15), .B(B_15), .C(C_15), .D(D_15), .E(E_15), .w_out(weight_2_15), .f_out(feature_2_15), .wf_en(wf_en_2_15), .opsum(psum_2_15));
	PEv2 # (.WIDTH(iWidth)) p_2_16(.clk(clk), .rst(rst), .in_en(wf_en_2_15), .ipsum(psum_3_16), .iconfig(iconfig_2), .weight(weight_2_15), .feature(feature_3_15), .config_load(config_load), .A(A_16), .B(B_16), .C(C_16), .D(D_16), .E(E_16), .w_out(weight_2_16), .f_out(feature_2_16), .wf_en(wf_en_2_16), .opsum(psum_2_16));
	PEv2 # (.WIDTH(iWidth)) p_2_17(.clk(clk), .rst(rst), .in_en(wf_en_2_16), .ipsum(psum_3_17), .iconfig(iconfig_2), .weight(weight_2_16), .feature(feature_3_16), .config_load(config_load), .A(A_17), .B(B_17), .C(C_17), .D(D_17), .E(E_17), .w_out(weight_2_17), .f_out(feature_2_17), .wf_en(wf_en_2_17), .opsum(psum_2_17));
	PEv2 # (.WIDTH(iWidth)) p_2_18(.clk(clk), .rst(rst), .in_en(wf_en_2_17), .ipsum(psum_3_18), .iconfig(iconfig_2), .weight(weight_2_17), .feature(feature_3_17), .config_load(config_load), .A(A_18), .B(B_18), .C(C_18), .D(D_18), .E(E_18), .w_out(weight_2_18), .f_out(feature_2_18), .wf_en(wf_en_2_18), .opsum(psum_2_18));
	PEv2 # (.WIDTH(iWidth)) p_2_19(.clk(clk), .rst(rst), .in_en(wf_en_2_18), .ipsum(psum_3_19), .iconfig(iconfig_2), .weight(weight_2_18), .feature(feature_3_18), .config_load(config_load), .A(A_19), .B(B_19), .C(C_19), .D(D_19), .E(E_19), .w_out(weight_2_19), .f_out(feature_2_19), .wf_en(wf_en_2_19), .opsum(psum_2_19));
	PEv2 # (.WIDTH(iWidth)) p_2_20(.clk(clk), .rst(rst), .in_en(wf_en_2_19), .ipsum(psum_3_20), .iconfig(iconfig_2), .weight(weight_2_19), .feature(feature_3_19), .config_load(config_load), .A(A_20), .B(B_20), .C(C_20), .D(D_20), .E(E_20), .w_out(weight_2_20), .f_out(feature_2_20), .wf_en(wf_en_2_20), .opsum(psum_2_20));
	PEv2 # (.WIDTH(iWidth)) p_2_21(.clk(clk), .rst(rst), .in_en(wf_en_2_20), .ipsum(psum_3_21), .iconfig(iconfig_2), .weight(weight_2_20), .feature(feature_3_20), .config_load(config_load), .A(A_21), .B(B_21), .C(C_21), .D(D_21), .E(E_21), .w_out(weight_2_21), .f_out(feature_2_21), .wf_en(wf_en_2_21), .opsum(psum_2_21));
	PEv2 # (.WIDTH(iWidth)) p_2_22(.clk(clk), .rst(rst), .in_en(wf_en_2_21), .ipsum(psum_3_22), .iconfig(iconfig_2), .weight(weight_2_21), .feature(feature_3_21), .config_load(config_load), .A(A_22), .B(B_22), .C(C_22), .D(D_22), .E(E_22), .w_out(weight_2_22), .f_out(feature_2_22), .wf_en(wf_en_2_22), .opsum(psum_2_22));
	PEv2 # (.WIDTH(iWidth)) p_2_23(.clk(clk), .rst(rst), .in_en(wf_en_2_22), .ipsum(psum_3_23), .iconfig(iconfig_2), .weight(weight_2_22), .feature(feature_3_22), .config_load(config_load), .A(A_23), .B(B_23), .C(C_23), .D(D_23), .E(E_23), .w_out(weight_2_23), .f_out(feature_2_23), .wf_en(wf_en_2_23), .opsum(psum_2_23));
	PEv2 # (.WIDTH(iWidth)) p_2_24(.clk(clk), .rst(rst), .in_en(wf_en_2_23), .ipsum(psum_3_24), .iconfig(iconfig_2), .weight(weight_2_23), .feature(feature_3_23), .config_load(config_load), .A(A_24), .B(B_24), .C(C_24), .D(D_24), .E(E_24), .w_out(weight_2_24), .f_out(feature_2_24), .wf_en(wf_en_2_24), .opsum(psum_2_24));
	PEv2 # (.WIDTH(iWidth)) p_2_25(.clk(clk), .rst(rst), .in_en(wf_en_2_24), .ipsum(psum_3_25), .iconfig(iconfig_2), .weight(weight_2_24), .feature(feature_3_24), .config_load(config_load), .A(A_25), .B(B_25), .C(C_25), .D(D_25), .E(E_25), .w_out(weight_2_25), .f_out(feature_2_25), .wf_en(wf_en_2_25), .opsum(psum_2_25));
	PEv2 # (.WIDTH(iWidth)) p_2_26(.clk(clk), .rst(rst), .in_en(wf_en_2_25), .ipsum(psum_3_26), .iconfig(iconfig_2), .weight(weight_2_25), .feature(feature_3_25), .config_load(config_load), .A(A_26), .B(B_26), .C(C_26), .D(D_26), .E(E_26), .w_out(weight_2_26), .f_out(feature_2_26), .wf_en(wf_en_2_26), .opsum(psum_2_26));
	PEv2 # (.WIDTH(iWidth)) p_2_27(.clk(clk), .rst(rst), .in_en(wf_en_2_26), .ipsum(psum_3_27), .iconfig(iconfig_2), .weight(weight_2_26), .feature(feature_3_26), .config_load(config_load), .A(A_27), .B(B_27), .C(C_27), .D(D_27), .E(E_27), .w_out(weight_2_27), .f_out(feature_2_27), .wf_en(wf_en_2_27), .opsum(psum_2_27));
	PEv2 # (.WIDTH(iWidth)) p_2_28(.clk(clk), .rst(rst), .in_en(wf_en_2_27), .ipsum(psum_3_28), .iconfig(iconfig_2), .weight(weight_2_27), .feature(feature_3_27), .config_load(config_load), .A(A_28), .B(B_28), .C(C_28), .D(D_28), .E(E_28), .w_out(weight_2_28), .f_out(feature_2_28), .wf_en(wf_en_2_28), .opsum(psum_2_28));
	PEv2 # (.WIDTH(iWidth)) p_2_29(.clk(clk), .rst(rst), .in_en(wf_en_2_28), .ipsum(psum_3_29), .iconfig(iconfig_2), .weight(weight_2_28), .feature(feature_3_28), .config_load(config_load), .A(A_29), .B(B_29), .C(C_29), .D(D_29), .E(E_29), .w_out(weight_2_29), .f_out(feature_2_29), .wf_en(wf_en_2_29), .opsum(psum_2_29));
	PEv2 # (.WIDTH(iWidth)) p_2_30(.clk(clk), .rst(rst), .in_en(wf_en_2_29), .ipsum(psum_3_30), .iconfig(iconfig_2), .weight(weight_2_29), .feature(feature_3_29), .config_load(config_load), .A(A_30), .B(B_30), .C(C_30), .D(D_30), .E(E_30), .w_out(weight_2_30), .f_out(feature_2_30), .wf_en(wf_en_2_30), .opsum(psum_2_30));
	PEv2 # (.WIDTH(iWidth)) p_2_31(.clk(clk), .rst(rst), .in_en(wf_en_2_30), .ipsum(psum_3_31), .iconfig(iconfig_2), .weight(weight_2_30), .feature(feature_3_30), .config_load(config_load), .A(A_31), .B(B_31), .C(C_31), .D(D_31), .E(E_31), .w_out(weight_2_31), .f_out(feature_2_31), .wf_en(wf_en_2_31), .opsum(psum_2_31));
	PEv2 # (.WIDTH(iWidth)) p_2_32(.clk(clk), .rst(rst), .in_en(wf_en_2_31), .ipsum(psum_3_32), .iconfig(iconfig_2), .weight(weight_2_31), .feature(feature_3_31), .config_load(config_load), .A(A_32), .B(B_32), .C(C_32), .D(D_32), .E(E_32), .w_out(weight_2_32), .f_out(feature_2_32), .wf_en(wf_en_2_32), .opsum(psum_2_32));
	PEv2 # (.WIDTH(iWidth)) p_3_1(.clk(clk), .rst(rst), .in_en(wf_en_3_0), .ipsum(psum_4_1), .iconfig(iconfig_3), .weight(weight_3_0), .feature(feature_4_0), .config_load(config_load), .A(A_1), .B(B_1), .C(C_1), .D(D_1), .E(E_1), .w_out(weight_3_1), .f_out(feature_3_1), .wf_en(wf_en_3_1), .opsum(psum_3_1));
	PEv2 # (.WIDTH(iWidth)) p_3_2(.clk(clk), .rst(rst), .in_en(wf_en_3_1), .ipsum(psum_4_2), .iconfig(iconfig_3), .weight(weight_3_1), .feature(feature_4_1), .config_load(config_load), .A(A_2), .B(B_2), .C(C_2), .D(D_2), .E(E_2), .w_out(weight_3_2), .f_out(feature_3_2), .wf_en(wf_en_3_2), .opsum(psum_3_2));
	PEv2 # (.WIDTH(iWidth)) p_3_3(.clk(clk), .rst(rst), .in_en(wf_en_3_2), .ipsum(psum_4_3), .iconfig(iconfig_3), .weight(weight_3_2), .feature(feature_4_2), .config_load(config_load), .A(A_3), .B(B_3), .C(C_3), .D(D_3), .E(E_3), .w_out(weight_3_3), .f_out(feature_3_3), .wf_en(wf_en_3_3), .opsum(psum_3_3));
	PEv2 # (.WIDTH(iWidth)) p_3_4(.clk(clk), .rst(rst), .in_en(wf_en_3_3), .ipsum(psum_4_4), .iconfig(iconfig_3), .weight(weight_3_3), .feature(feature_4_3), .config_load(config_load), .A(A_4), .B(B_4), .C(C_4), .D(D_4), .E(E_4), .w_out(weight_3_4), .f_out(feature_3_4), .wf_en(wf_en_3_4), .opsum(psum_3_4));
	PEv2 # (.WIDTH(iWidth)) p_3_5(.clk(clk), .rst(rst), .in_en(wf_en_3_4), .ipsum(psum_4_5), .iconfig(iconfig_3), .weight(weight_3_4), .feature(feature_4_4), .config_load(config_load), .A(A_5), .B(B_5), .C(C_5), .D(D_5), .E(E_5), .w_out(weight_3_5), .f_out(feature_3_5), .wf_en(wf_en_3_5), .opsum(psum_3_5));
	PEv2 # (.WIDTH(iWidth)) p_3_6(.clk(clk), .rst(rst), .in_en(wf_en_3_5), .ipsum(psum_4_6), .iconfig(iconfig_3), .weight(weight_3_5), .feature(feature_4_5), .config_load(config_load), .A(A_6), .B(B_6), .C(C_6), .D(D_6), .E(E_6), .w_out(weight_3_6), .f_out(feature_3_6), .wf_en(wf_en_3_6), .opsum(psum_3_6));
	PEv2 # (.WIDTH(iWidth)) p_3_7(.clk(clk), .rst(rst), .in_en(wf_en_3_6), .ipsum(psum_4_7), .iconfig(iconfig_3), .weight(weight_3_6), .feature(feature_4_6), .config_load(config_load), .A(A_7), .B(B_7), .C(C_7), .D(D_7), .E(E_7), .w_out(weight_3_7), .f_out(feature_3_7), .wf_en(wf_en_3_7), .opsum(psum_3_7));
	PEv2 # (.WIDTH(iWidth)) p_3_8(.clk(clk), .rst(rst), .in_en(wf_en_3_7), .ipsum(psum_4_8), .iconfig(iconfig_3), .weight(weight_3_7), .feature(feature_4_7), .config_load(config_load), .A(A_8), .B(B_8), .C(C_8), .D(D_8), .E(E_8), .w_out(weight_3_8), .f_out(feature_3_8), .wf_en(wf_en_3_8), .opsum(psum_3_8));
	PEv2 # (.WIDTH(iWidth)) p_3_9(.clk(clk), .rst(rst), .in_en(wf_en_3_8), .ipsum(psum_4_9), .iconfig(iconfig_3), .weight(weight_3_8), .feature(feature_4_8), .config_load(config_load), .A(A_9), .B(B_9), .C(C_9), .D(D_9), .E(E_9), .w_out(weight_3_9), .f_out(feature_3_9), .wf_en(wf_en_3_9), .opsum(psum_3_9));
	PEv2 # (.WIDTH(iWidth)) p_3_10(.clk(clk), .rst(rst), .in_en(wf_en_3_9), .ipsum(psum_4_10), .iconfig(iconfig_3), .weight(weight_3_9), .feature(feature_4_9), .config_load(config_load), .A(A_10), .B(B_10), .C(C_10), .D(D_10), .E(E_10), .w_out(weight_3_10), .f_out(feature_3_10), .wf_en(wf_en_3_10), .opsum(psum_3_10));
	PEv2 # (.WIDTH(iWidth)) p_3_11(.clk(clk), .rst(rst), .in_en(wf_en_3_10), .ipsum(psum_4_11), .iconfig(iconfig_3), .weight(weight_3_10), .feature(feature_4_10), .config_load(config_load), .A(A_11), .B(B_11), .C(C_11), .D(D_11), .E(E_11), .w_out(weight_3_11), .f_out(feature_3_11), .wf_en(wf_en_3_11), .opsum(psum_3_11));
	PEv2 # (.WIDTH(iWidth)) p_3_12(.clk(clk), .rst(rst), .in_en(wf_en_3_11), .ipsum(psum_4_12), .iconfig(iconfig_3), .weight(weight_3_11), .feature(feature_4_11), .config_load(config_load), .A(A_12), .B(B_12), .C(C_12), .D(D_12), .E(E_12), .w_out(weight_3_12), .f_out(feature_3_12), .wf_en(wf_en_3_12), .opsum(psum_3_12));
	PEv2 # (.WIDTH(iWidth)) p_3_13(.clk(clk), .rst(rst), .in_en(wf_en_3_12), .ipsum(psum_4_13), .iconfig(iconfig_3), .weight(weight_3_12), .feature(feature_4_12), .config_load(config_load), .A(A_13), .B(B_13), .C(C_13), .D(D_13), .E(E_13), .w_out(weight_3_13), .f_out(feature_3_13), .wf_en(wf_en_3_13), .opsum(psum_3_13));
	PEv2 # (.WIDTH(iWidth)) p_3_14(.clk(clk), .rst(rst), .in_en(wf_en_3_13), .ipsum(psum_4_14), .iconfig(iconfig_3), .weight(weight_3_13), .feature(feature_4_13), .config_load(config_load), .A(A_14), .B(B_14), .C(C_14), .D(D_14), .E(E_14), .w_out(weight_3_14), .f_out(feature_3_14), .wf_en(wf_en_3_14), .opsum(psum_3_14));
	PEv2 # (.WIDTH(iWidth)) p_3_15(.clk(clk), .rst(rst), .in_en(wf_en_3_14), .ipsum(psum_4_15), .iconfig(iconfig_3), .weight(weight_3_14), .feature(feature_4_14), .config_load(config_load), .A(A_15), .B(B_15), .C(C_15), .D(D_15), .E(E_15), .w_out(weight_3_15), .f_out(feature_3_15), .wf_en(wf_en_3_15), .opsum(psum_3_15));
	PEv2 # (.WIDTH(iWidth)) p_3_16(.clk(clk), .rst(rst), .in_en(wf_en_3_15), .ipsum(psum_4_16), .iconfig(iconfig_3), .weight(weight_3_15), .feature(feature_4_15), .config_load(config_load), .A(A_16), .B(B_16), .C(C_16), .D(D_16), .E(E_16), .w_out(weight_3_16), .f_out(feature_3_16), .wf_en(wf_en_3_16), .opsum(psum_3_16));
	PEv2 # (.WIDTH(iWidth)) p_3_17(.clk(clk), .rst(rst), .in_en(wf_en_3_16), .ipsum(psum_4_17), .iconfig(iconfig_3), .weight(weight_3_16), .feature(feature_4_16), .config_load(config_load), .A(A_17), .B(B_17), .C(C_17), .D(D_17), .E(E_17), .w_out(weight_3_17), .f_out(feature_3_17), .wf_en(wf_en_3_17), .opsum(psum_3_17));
	PEv2 # (.WIDTH(iWidth)) p_3_18(.clk(clk), .rst(rst), .in_en(wf_en_3_17), .ipsum(psum_4_18), .iconfig(iconfig_3), .weight(weight_3_17), .feature(feature_4_17), .config_load(config_load), .A(A_18), .B(B_18), .C(C_18), .D(D_18), .E(E_18), .w_out(weight_3_18), .f_out(feature_3_18), .wf_en(wf_en_3_18), .opsum(psum_3_18));
	PEv2 # (.WIDTH(iWidth)) p_3_19(.clk(clk), .rst(rst), .in_en(wf_en_3_18), .ipsum(psum_4_19), .iconfig(iconfig_3), .weight(weight_3_18), .feature(feature_4_18), .config_load(config_load), .A(A_19), .B(B_19), .C(C_19), .D(D_19), .E(E_19), .w_out(weight_3_19), .f_out(feature_3_19), .wf_en(wf_en_3_19), .opsum(psum_3_19));
	PEv2 # (.WIDTH(iWidth)) p_3_20(.clk(clk), .rst(rst), .in_en(wf_en_3_19), .ipsum(psum_4_20), .iconfig(iconfig_3), .weight(weight_3_19), .feature(feature_4_19), .config_load(config_load), .A(A_20), .B(B_20), .C(C_20), .D(D_20), .E(E_20), .w_out(weight_3_20), .f_out(feature_3_20), .wf_en(wf_en_3_20), .opsum(psum_3_20));
	PEv2 # (.WIDTH(iWidth)) p_3_21(.clk(clk), .rst(rst), .in_en(wf_en_3_20), .ipsum(psum_4_21), .iconfig(iconfig_3), .weight(weight_3_20), .feature(feature_4_20), .config_load(config_load), .A(A_21), .B(B_21), .C(C_21), .D(D_21), .E(E_21), .w_out(weight_3_21), .f_out(feature_3_21), .wf_en(wf_en_3_21), .opsum(psum_3_21));
	PEv2 # (.WIDTH(iWidth)) p_3_22(.clk(clk), .rst(rst), .in_en(wf_en_3_21), .ipsum(psum_4_22), .iconfig(iconfig_3), .weight(weight_3_21), .feature(feature_4_21), .config_load(config_load), .A(A_22), .B(B_22), .C(C_22), .D(D_22), .E(E_22), .w_out(weight_3_22), .f_out(feature_3_22), .wf_en(wf_en_3_22), .opsum(psum_3_22));
	PEv2 # (.WIDTH(iWidth)) p_3_23(.clk(clk), .rst(rst), .in_en(wf_en_3_22), .ipsum(psum_4_23), .iconfig(iconfig_3), .weight(weight_3_22), .feature(feature_4_22), .config_load(config_load), .A(A_23), .B(B_23), .C(C_23), .D(D_23), .E(E_23), .w_out(weight_3_23), .f_out(feature_3_23), .wf_en(wf_en_3_23), .opsum(psum_3_23));
	PEv2 # (.WIDTH(iWidth)) p_3_24(.clk(clk), .rst(rst), .in_en(wf_en_3_23), .ipsum(psum_4_24), .iconfig(iconfig_3), .weight(weight_3_23), .feature(feature_4_23), .config_load(config_load), .A(A_24), .B(B_24), .C(C_24), .D(D_24), .E(E_24), .w_out(weight_3_24), .f_out(feature_3_24), .wf_en(wf_en_3_24), .opsum(psum_3_24));
	PEv2 # (.WIDTH(iWidth)) p_3_25(.clk(clk), .rst(rst), .in_en(wf_en_3_24), .ipsum(psum_4_25), .iconfig(iconfig_3), .weight(weight_3_24), .feature(feature_4_24), .config_load(config_load), .A(A_25), .B(B_25), .C(C_25), .D(D_25), .E(E_25), .w_out(weight_3_25), .f_out(feature_3_25), .wf_en(wf_en_3_25), .opsum(psum_3_25));
	PEv2 # (.WIDTH(iWidth)) p_3_26(.clk(clk), .rst(rst), .in_en(wf_en_3_25), .ipsum(psum_4_26), .iconfig(iconfig_3), .weight(weight_3_25), .feature(feature_4_25), .config_load(config_load), .A(A_26), .B(B_26), .C(C_26), .D(D_26), .E(E_26), .w_out(weight_3_26), .f_out(feature_3_26), .wf_en(wf_en_3_26), .opsum(psum_3_26));
	PEv2 # (.WIDTH(iWidth)) p_3_27(.clk(clk), .rst(rst), .in_en(wf_en_3_26), .ipsum(psum_4_27), .iconfig(iconfig_3), .weight(weight_3_26), .feature(feature_4_26), .config_load(config_load), .A(A_27), .B(B_27), .C(C_27), .D(D_27), .E(E_27), .w_out(weight_3_27), .f_out(feature_3_27), .wf_en(wf_en_3_27), .opsum(psum_3_27));
	PEv2 # (.WIDTH(iWidth)) p_3_28(.clk(clk), .rst(rst), .in_en(wf_en_3_27), .ipsum(psum_4_28), .iconfig(iconfig_3), .weight(weight_3_27), .feature(feature_4_27), .config_load(config_load), .A(A_28), .B(B_28), .C(C_28), .D(D_28), .E(E_28), .w_out(weight_3_28), .f_out(feature_3_28), .wf_en(wf_en_3_28), .opsum(psum_3_28));
	PEv2 # (.WIDTH(iWidth)) p_3_29(.clk(clk), .rst(rst), .in_en(wf_en_3_28), .ipsum(psum_4_29), .iconfig(iconfig_3), .weight(weight_3_28), .feature(feature_4_28), .config_load(config_load), .A(A_29), .B(B_29), .C(C_29), .D(D_29), .E(E_29), .w_out(weight_3_29), .f_out(feature_3_29), .wf_en(wf_en_3_29), .opsum(psum_3_29));
	PEv2 # (.WIDTH(iWidth)) p_3_30(.clk(clk), .rst(rst), .in_en(wf_en_3_29), .ipsum(psum_4_30), .iconfig(iconfig_3), .weight(weight_3_29), .feature(feature_4_29), .config_load(config_load), .A(A_30), .B(B_30), .C(C_30), .D(D_30), .E(E_30), .w_out(weight_3_30), .f_out(feature_3_30), .wf_en(wf_en_3_30), .opsum(psum_3_30));
	PEv2 # (.WIDTH(iWidth)) p_3_31(.clk(clk), .rst(rst), .in_en(wf_en_3_30), .ipsum(psum_4_31), .iconfig(iconfig_3), .weight(weight_3_30), .feature(feature_4_30), .config_load(config_load), .A(A_31), .B(B_31), .C(C_31), .D(D_31), .E(E_31), .w_out(weight_3_31), .f_out(feature_3_31), .wf_en(wf_en_3_31), .opsum(psum_3_31));
	PEv2 # (.WIDTH(iWidth)) p_3_32(.clk(clk), .rst(rst), .in_en(wf_en_3_31), .ipsum(psum_4_32), .iconfig(iconfig_3), .weight(weight_3_31), .feature(feature_4_31), .config_load(config_load), .A(A_32), .B(B_32), .C(C_32), .D(D_32), .E(E_32), .w_out(weight_3_32), .f_out(feature_3_32), .wf_en(wf_en_3_32), .opsum(psum_3_32));

	AC # (.IN_WIDTH(oWidth), .ACC_WIDTH(oWidth)) ac_1(.clk(clk), .rst(rst), .in_en(G_1), .ipsum(psum_1_1), .F(F_1), .data_out(dout_1));
	AC # (.IN_WIDTH(oWidth), .ACC_WIDTH(oWidth)) ac_2(.clk(clk), .rst(rst), .in_en(G_2), .ipsum(psum_1_2), .F(F_2), .data_out(dout_2));
	AC # (.IN_WIDTH(oWidth), .ACC_WIDTH(oWidth)) ac_3(.clk(clk), .rst(rst), .in_en(G_3), .ipsum(psum_1_3), .F(F_3), .data_out(dout_3));
	AC # (.IN_WIDTH(oWidth), .ACC_WIDTH(oWidth)) ac_4(.clk(clk), .rst(rst), .in_en(G_4), .ipsum(psum_1_4), .F(F_4), .data_out(dout_4));
	AC # (.IN_WIDTH(oWidth), .ACC_WIDTH(oWidth)) ac_5(.clk(clk), .rst(rst), .in_en(G_5), .ipsum(psum_1_5), .F(F_5), .data_out(dout_5));
	AC # (.IN_WIDTH(oWidth), .ACC_WIDTH(oWidth)) ac_6(.clk(clk), .rst(rst), .in_en(G_6), .ipsum(psum_1_6), .F(F_6), .data_out(dout_6));
	AC # (.IN_WIDTH(oWidth), .ACC_WIDTH(oWidth)) ac_7(.clk(clk), .rst(rst), .in_en(G_7), .ipsum(psum_1_7), .F(F_7), .data_out(dout_7));
	AC # (.IN_WIDTH(oWidth), .ACC_WIDTH(oWidth)) ac_8(.clk(clk), .rst(rst), .in_en(G_8), .ipsum(psum_1_8), .F(F_8), .data_out(dout_8));
	AC # (.IN_WIDTH(oWidth), .ACC_WIDTH(oWidth)) ac_9(.clk(clk), .rst(rst), .in_en(G_9), .ipsum(psum_1_9), .F(F_9), .data_out(dout_9));
	AC # (.IN_WIDTH(oWidth), .ACC_WIDTH(oWidth)) ac_10(.clk(clk), .rst(rst), .in_en(G_10), .ipsum(psum_1_10), .F(F_10), .data_out(dout_10));
	AC # (.IN_WIDTH(oWidth), .ACC_WIDTH(oWidth)) ac_11(.clk(clk), .rst(rst), .in_en(G_11), .ipsum(psum_1_11), .F(F_11), .data_out(dout_11));
	AC # (.IN_WIDTH(oWidth), .ACC_WIDTH(oWidth)) ac_12(.clk(clk), .rst(rst), .in_en(G_12), .ipsum(psum_1_12), .F(F_12), .data_out(dout_12));
	AC # (.IN_WIDTH(oWidth), .ACC_WIDTH(oWidth)) ac_13(.clk(clk), .rst(rst), .in_en(G_13), .ipsum(psum_1_13), .F(F_13), .data_out(dout_13));
	AC # (.IN_WIDTH(oWidth), .ACC_WIDTH(oWidth)) ac_14(.clk(clk), .rst(rst), .in_en(G_14), .ipsum(psum_1_14), .F(F_14), .data_out(dout_14));
	AC # (.IN_WIDTH(oWidth), .ACC_WIDTH(oWidth)) ac_15(.clk(clk), .rst(rst), .in_en(G_15), .ipsum(psum_1_15), .F(F_15), .data_out(dout_15));
	AC # (.IN_WIDTH(oWidth), .ACC_WIDTH(oWidth)) ac_16(.clk(clk), .rst(rst), .in_en(G_16), .ipsum(psum_1_16), .F(F_16), .data_out(dout_16));
	AC # (.IN_WIDTH(oWidth), .ACC_WIDTH(oWidth)) ac_17(.clk(clk), .rst(rst), .in_en(G_17), .ipsum(psum_1_17), .F(F_17), .data_out(dout_17));
	AC # (.IN_WIDTH(oWidth), .ACC_WIDTH(oWidth)) ac_18(.clk(clk), .rst(rst), .in_en(G_18), .ipsum(psum_1_18), .F(F_18), .data_out(dout_18));
	AC # (.IN_WIDTH(oWidth), .ACC_WIDTH(oWidth)) ac_19(.clk(clk), .rst(rst), .in_en(G_19), .ipsum(psum_1_19), .F(F_19), .data_out(dout_19));
	AC # (.IN_WIDTH(oWidth), .ACC_WIDTH(oWidth)) ac_20(.clk(clk), .rst(rst), .in_en(G_20), .ipsum(psum_1_20), .F(F_20), .data_out(dout_20));
	AC # (.IN_WIDTH(oWidth), .ACC_WIDTH(oWidth)) ac_21(.clk(clk), .rst(rst), .in_en(G_21), .ipsum(psum_1_21), .F(F_21), .data_out(dout_21));
	AC # (.IN_WIDTH(oWidth), .ACC_WIDTH(oWidth)) ac_22(.clk(clk), .rst(rst), .in_en(G_22), .ipsum(psum_1_22), .F(F_22), .data_out(dout_22));
	AC # (.IN_WIDTH(oWidth), .ACC_WIDTH(oWidth)) ac_23(.clk(clk), .rst(rst), .in_en(G_23), .ipsum(psum_1_23), .F(F_23), .data_out(dout_23));
	AC # (.IN_WIDTH(oWidth), .ACC_WIDTH(oWidth)) ac_24(.clk(clk), .rst(rst), .in_en(G_24), .ipsum(psum_1_24), .F(F_24), .data_out(dout_24));
	AC # (.IN_WIDTH(oWidth), .ACC_WIDTH(oWidth)) ac_25(.clk(clk), .rst(rst), .in_en(G_25), .ipsum(psum_1_25), .F(F_25), .data_out(dout_25));
	AC # (.IN_WIDTH(oWidth), .ACC_WIDTH(oWidth)) ac_26(.clk(clk), .rst(rst), .in_en(G_26), .ipsum(psum_1_26), .F(F_26), .data_out(dout_26));
	AC # (.IN_WIDTH(oWidth), .ACC_WIDTH(oWidth)) ac_27(.clk(clk), .rst(rst), .in_en(G_27), .ipsum(psum_1_27), .F(F_27), .data_out(dout_27));
	AC # (.IN_WIDTH(oWidth), .ACC_WIDTH(oWidth)) ac_28(.clk(clk), .rst(rst), .in_en(G_28), .ipsum(psum_1_28), .F(F_28), .data_out(dout_28));
	AC # (.IN_WIDTH(oWidth), .ACC_WIDTH(oWidth)) ac_29(.clk(clk), .rst(rst), .in_en(G_29), .ipsum(psum_1_29), .F(F_29), .data_out(dout_29));
	AC # (.IN_WIDTH(oWidth), .ACC_WIDTH(oWidth)) ac_30(.clk(clk), .rst(rst), .in_en(G_30), .ipsum(psum_1_30), .F(F_30), .data_out(dout_30));
	AC # (.IN_WIDTH(oWidth), .ACC_WIDTH(oWidth)) ac_31(.clk(clk), .rst(rst), .in_en(G_31), .ipsum(psum_1_31), .F(F_31), .data_out(dout_31));
	AC # (.IN_WIDTH(oWidth), .ACC_WIDTH(oWidth)) ac_32(.clk(clk), .rst(rst), .in_en(G_32), .ipsum(psum_1_32), .F(F_32), .data_out(dout_32));
endmodule
